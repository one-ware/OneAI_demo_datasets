library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.numeric_std.all;
use work.CNN_Config_Package.all;

PACKAGE CNN_Data_Package is
  CONSTANT Layer_1_Columns    : NATURAL := 128;
  CONSTANT Layer_1_Rows       : NATURAL := 128;
  CONSTANT Layer_1_Strides    : NATURAL := 1;
  CONSTANT Layer_1_Activation : Activation_T := relu;
  CONSTANT Layer_1_Padding    : Padding_T := same;
  CONSTANT Layer_1_Values     : NATURAL := 1;
  CONSTANT Layer_1_Filter_X   : NATURAL := 3;
  CONSTANT Layer_1_Filter_Y   : NATURAL := 3;
  CONSTANT Layer_1_Filters    : NATURAL := 8;
  CONSTANT Layer_1_Inputs     : NATURAL := 10;
  CONSTANT Layer_1_Out_Offset : INTEGER := 3;
  CONSTANT Layer_1_Offset     : INTEGER := 1;
  CONSTANT Layer_1 : CNN_Weights_T(0 to Layer_1_Filters-1, 0 to Layer_1_Inputs-1) :=
  (
    (-33, -39, -41, -39, -32, -39, -10, -2, -37, 0),
    (-49, -27, -16, 13, 68, -25, -34, 8, -49, -1),
    (7, 21, 6, -11, 1, 20, -7, 33, -2, -1),
    (-77, -81, -33, -5, -20, -15, 21, 45, 18, 1),
    (64, -40, -54, 13, 2, 1, 31, 15, -10, -7),
    (39, 23, 27, 18, -8, -32, -14, -39, -59, -1),
    (23, 44, -11, 6, 24, 21, -7, -10, 10, -7),
    (11, -18, 28, -1, 20, 18, 4, -15, 49, -5)
  );
  ----------------
  CONSTANT Pooling_1_Columns      : NATURAL := 128;
  CONSTANT Pooling_1_Rows         : NATURAL := 128;
  CONSTANT Pooling_1_Values       : NATURAL := 8;
  CONSTANT Pooling_1_Filter_X     : NATURAL := 2;
  CONSTANT Pooling_1_Filter_Y     : NATURAL := 2;
  CONSTANT Pooling_1_Strides      : NATURAL := 2;
  CONSTANT Pooling_1_Padding      : Padding_T := valid;
  ----------------
  CONSTANT Layer_2_Columns    : NATURAL := 64;
  CONSTANT Layer_2_Rows       : NATURAL := 64;
  CONSTANT Layer_2_Strides    : NATURAL := 2;
  CONSTANT Layer_2_Activation : Activation_T := relu;
  CONSTANT Layer_2_Padding    : Padding_T := same;
  CONSTANT Layer_2_Values     : NATURAL := 8;
  CONSTANT Layer_2_Filter_X   : NATURAL := 3;
  CONSTANT Layer_2_Filter_Y   : NATURAL := 3;
  CONSTANT Layer_2_Filters    : NATURAL := 12;
  CONSTANT Layer_2_Inputs     : NATURAL := 73;
  CONSTANT Layer_2_Out_Offset : INTEGER := 4;
  CONSTANT Layer_2_Offset     : INTEGER := 1;
  CONSTANT Layer_2 : CNN_Weights_T(0 to Layer_2_Filters-1, 0 to Layer_2_Inputs-1) :=
  (
    (1, -3, -2, 5, 5, 2, 9, -3, 1, 7, -6, 16, 15, -2, 15, -16, -15, -19, -23, -18, 3, 10, 1, -17, 5, 16, 21, -19, 22, 3, 20, 17, 6, 13, 3, -12, 14, 14, 6, -12, 13, -38, -7, 0, -28, 30, -7, -30, -6, 19, 6, -3, 24, -4, 21, 0, 15, -3, -10, -26, 10, 14, -9, -1, 14, -32, -7, 19, -21, -10, -6, -5, -1),
    (-1, 10, -26, 26, 18, -7, -7, -12, 5, -14, -25, 14, 2, -17, -19, -25, -3, -22, -2, -15, -13, 36, -15, -22, 13, 20, 20, 3, 33, 22, 12, 24, -8, 2, -3, 5, 15, -25, 6, 12, 13, -1, -9, -9, 2, -27, -15, -13, 9, 15, 16, -1, -5, 14, 11, 13, -2, 24, -1, 14, 6, -7, 21, -6, -2, 15, -2, 16, 17, -19, 8, -3, -4),
    (6, 23, -6, 26, -29, -46, -12, 17, -5, 31, 23, -5, -26, -94, 1, 19, -12, 13, 17, -11, -14, -38, -6, 9, -17, 29, -6, 1, -7, -82, 6, -4, -1, 33, -8, 1, -10, -90, 5, 9, -15, 16, 19, -12, 9, -50, 2, 13, -8, 4, -8, -11, -7, -38, 11, 11, 12, -3, -4, 5, -5, -50, 3, 6, 9, -6, 17, 14, 17, -25, -2, 12, 0),
    (-12, 1, 15, -15, 18, 14, 18, 2, 13, 7, 1, -24, -5, 2, 8, 12, -14, 20, 11, -12, 7, -12, -2, 4, 3, 14, -4, -16, 31, 1, 9, 6, 2, 15, 0, -17, 6, -5, 22, 6, 18, 26, -2, -9, 11, 2, -1, 17, 7, 14, -4, -10, 6, 8, 10, 6, 10, 24, 9, -12, 6, -6, 8, -14, -8, 27, -6, -5, 11, 10, -2, -11, -2),
    (-14, 11, 10, -1, 5, 10, 0, 18, -16, 13, 10, 16, 1, 15, 20, 21, -12, -12, 22, 23, -6, 18, 22, 13, 13, 1, 3, 21, -18, 15, -13, -6, -7, -17, 4, 42, -20, 18, -4, -9, 6, -11, 16, 48, -13, 18, 9, 14, -1, -24, -5, 19, 7, -14, -16, -7, 1, -68, -22, 19, -9, 6, -31, -27, 5, -42, -20, 27, -20, 4, -15, -15, -6),
    (-8, 13, 6, -28, 22, 5, 1, 4, 8, -46, -29, -28, 7, -15, -16, -22, 1, 25, -6, -11, -12, -14, 4, 32, -7, 22, -25, -29, 26, 2, 2, -18, -1, -94, -10, -28, 6, -11, -18, -6, -1, 41, 17, -16, 1, -10, 14, 19, -14, 1, -14, -15, 5, 20, -2, -25, 1, -35, 10, -22, 0, -14, -8, 3, -17, 26, 15, -3, 11, -13, 6, 18, 0),
    (-17, 18, 15, -2, 12, 18, 14, 20, -14, 13, 8, -65, 11, 15, 2, 2, 13, -35, -19, -75, -14, -1, -5, -16, -17, 13, 6, 21, 21, 34, 14, 8, 1, 5, -8, -49, 5, 3, -10, -18, -10, -91, -14, -5, -4, 2, -15, -6, -13, -3, -27, 21, -17, 22, -14, -17, 7, -52, -8, 14, -23, 13, -6, -17, -6, -111, 13, 14, -8, -89, 9, 15, 0),
    (-1, 2, 15, -31, -6, -29, 12, 19, -5, 26, 13, -18, 22, -30, 13, -2, -6, 15, -22, 14, 23, -2, 0, -15, -13, 18, 2, -45, 4, -30, 5, 4, 15, 52, 15, -27, 22, -36, 17, 11, 9, 45, -1, -1, 24, -24, 5, -9, 7, -7, -9, -53, -19, -31, -18, -7, -11, 49, 0, -18, 4, -17, 19, 2, 16, 28, 8, -4, 10, -18, 17, 5, -6),
    (-16, 10, -17, 14, -4, -2, -29, -17, -6, 29, -9, 24, 5, 16, -2, 5, 17, 50, 2, 15, -8, -19, -14, -25, 0, 30, 4, 15, -20, 48, -19, -3, -7, 24, 5, 38, 0, 26, 8, -2, 0, 39, -6, -15, 10, -9, -7, -19, 17, 18, 15, 18, -17, 42, 5, 2, 2, 20, -1, 12, -1, 20, 4, -12, -12, 13, -44, -36, 14, 1, -8, -40, 0),
    (-9, -52, -20, -13, -5, 41, -26, -18, -10, 18, -10, 10, -19, -46, -15, 2, 1, -4, 2, 19, -8, -6, -3, -6, 14, -61, 1, 12, -2, -30, -5, -8, 17, 18, 27, -3, -14, -4, -3, 10, 12, 4, 11, 11, 9, 29, -7, 8, -2, -7, -1, 5, -9, -22, -11, 18, -6, 35, 11, -3, -11, -7, 22, 3, -15, 18, -8, -8, 12, 23, 12, 6, 2),
    (7, 9, 10, 28, -10, -12, -5, -7, -3, -7, 5, 14, 13, -2, -8, 8, 10, -24, 8, 10, -6, -2, -6, 6, 12, -10, 6, 9, -10, -5, 13, 11, -17, -8, 3, 16, -2, 10, 13, 4, 8, -24, 17, 16, -23, 10, -1, -2, 12, -6, -3, 17, 10, -1, 17, 11, 16, -26, -4, 22, -7, 2, 6, 14, -17, -37, 14, 15, -18, -6, -8, 23, -1),
    (7, 39, 8, -1, -15, -8, -12, 1, 4, 16, 1, -4, -10, -10, 9, 6, 10, -14, 2, -22, -19, 6, 15, 8, 0, 49, 15, -4, -16, -5, 15, 2, 10, 46, 11, -6, -8, 13, 4, 6, -1, 5, 13, 7, -15, 11, 19, 7, -10, 46, -7, -10, -16, -4, -10, 1, 8, 28, -4, 5, -11, 33, 0, 6, -15, 16, -2, -4, -12, 31, 5, -12, -3)
  );
  ----------------
  CONSTANT Layer_3_Columns    : NATURAL := 32;
  CONSTANT Layer_3_Rows       : NATURAL := 32;
  CONSTANT Layer_3_Strides    : NATURAL := 2;
  CONSTANT Layer_3_Activation : Activation_T := relu;
  CONSTANT Layer_3_Padding    : Padding_T := same;
  CONSTANT Layer_3_Values     : NATURAL := 12;
  CONSTANT Layer_3_Filter_X   : NATURAL := 3;
  CONSTANT Layer_3_Filter_Y   : NATURAL := 3;
  CONSTANT Layer_3_Filters    : NATURAL := 16;
  CONSTANT Layer_3_Inputs     : NATURAL := 109;
  CONSTANT Layer_3_Out_Offset : INTEGER := 5;
  CONSTANT Layer_3_Offset     : INTEGER := 1;
  CONSTANT Layer_3 : CNN_Weights_T(0 to Layer_3_Filters-1, 0 to Layer_3_Inputs-1) :=
  (
    (-19, 13, 0, -25, 14, 13, 9, -13, 22, 18, -14, -15, -16, 18, -21, -9, 18, 13, -3, -22, 12, 2, -11, -25, 6, -1, -14, -10, 10, 13, -13, -15, 1, 3, -16, -3, -45, -2, 10, -7, -80, -6, -6, -8, -26, 4, 3, -5, -33, 14, 5, -14, -55, -13, -18, 14, -30, -16, 0, -26, -9, 10, 9, -10, -14, 1, -6, 17, -14, -15, -3, -31, -2, 2, 2, 27, -6, 6, 5, 12, 7, -6, 17, 3, -10, 17, 19, 20, 0, -9, -13, 14, -6, 6, 21, 21, -15, 22, 22, 0, 10, -24, -6, 11, -10, -3, 18, 14, 4),
    (-1, 5, -7, 3, 3, -5, -4, 2, 5, -4, -8, 3, 6, 0, -16, 13, 9, 7, -3, 3, 13, -2, 4, -2, 6, -10, -2, 0, 13, 9, 4, 2, -1, 2, 20, 20, -5, 8, -18, 9, 4, 2, -2, -3, 23, 1, 2, 3, -7, 2, -11, 9, 22, -17, 0, -2, 14, -1, 1, 12, -6, -4, 10, 14, 17, 6, -10, -9, -10, 12, 25, 16, -7, 5, -6, -7, 10, -3, -12, 4, -4, 6, -14, 6, -5, -2, -16, -2, 10, -15, -7, 1, 16, 2, 14, 3, -1, -7, 3, 5, 6, -2, -2, 1, 5, -5, 12, 5, -3),
    (-43, 12, -15, 0, 14, -53, -27, -14, -6, -26, 8, -6, -36, 4, 12, 6, -13, -11, 0, -14, 2, -3, 6, -15, 1, -15, 7, 3, -3, 15, 4, -10, 1, 18, 12, 18, -56, -26, 14, -22, -5, -12, -2, -34, -37, 14, 10, -9, 7, -34, 15, 3, -31, -15, 33, -20, -16, 8, 10, 13, 8, -31, 8, 8, -2, 17, 14, -9, -1, 14, 6, 21, 9, -19, 19, 3, -14, 2, 9, 2, -4, 18, 10, -2, 24, -26, 10, 15, -13, 17, 22, -2, -8, 19, -6, 11, 10, -12, 10, 10, -2, 2, -9, -10, -7, 0, -14, 6, 0),
    (10, -10, -17, -13, -32, 14, 8, 16, -24, -9, -9, -1, 17, -7, 8, -23, -45, 7, -15, -35, -38, 0, -13, -17, -2, -14, 14, -2, -69, -13, 7, -22, 22, -5, -8, -2, -7, 10, -16, -19, -15, -17, 13, 14, -27, -28, -15, -41, -22, -3, 15, -8, -43, -3, 20, -28, 21, 4, -10, -8, 2, -8, 4, 11, -43, 12, 24, -11, 4, 10, 16, 3, 20, -6, 7, -13, -6, -25, 13, -14, 12, -10, 5, -9, 28, -4, 20, 9, -13, 16, 54, -18, 15, 11, 14, -5, 26, -8, 18, 22, -2, 31, 28, -2, 2, 14, -1, 14, 0),
    (3, -4, -10, -3, 5, 21, 23, 10, -8, 14, 8, 10, 14, -11, -4, -1, 2, 9, 7, 7, -24, 10, -5, 21, -6, -2, 2, 10, 3, -13, -11, 7, -21, -10, 7, 0, 10, -40, 2, -4, -16, 24, 31, -6, 24, 10, 0, 6, 22, -52, -2, 0, -10, 31, 29, -2, 13, 20, -10, -1, 13, -4, -18, 7, -2, 13, -8, -1, -22, 13, -15, -2, 5, -15, 6, 1, -17, 12, 17, -10, 19, 12, 13, -8, 16, -26, 0, 6, -24, 31, 30, -15, 26, 32, -1, 9, 2, -21, -26, -11, -5, 21, 19, -12, 11, 18, 10, 5, -19),
    (13, -12, 13, 16, -9, 9, 31, 8, -6, 9, 10, 1, 7, -15, -5, 11, 1, -2, 28, -8, 0, 18, 16, 2, -4, -2, -15, -3, 2, -16, 12, -22, 4, 18, -6, -4, 20, 7, 5, 10, -1, -1, -12, 22, -17, -1, -2, 0, 6, 1, -11, 18, -4, -38, -15, 10, 2, 0, 13, -4, 2, -7, -11, -3, 7, -26, -5, -14, 24, 4, 1, -18, 2, 15, -7, 5, 12, 2, -13, 31, -30, -23, 1, 0, -18, 25, 9, 1, 10, -28, -42, 19, -26, -23, 9, 14, -6, 10, 3, -13, 9, -52, -25, 3, -13, -14, -10, -6, 1),
    (-9, -29, 24, 14, -14, 12, 27, 5, 7, 4, 23, -5, 10, -50, 29, 1, -14, 27, 45, 2, -10, 43, 10, 24, -2, -30, -11, 2, -5, 0, 37, -9, -22, 44, -3, 10, 11, -48, 23, -2, -3, -9, 25, 8, 23, -6, 10, 14, 3, -81, -26, 2, -7, -2, 28, -34, -14, 9, 15, 6, -2, -48, -2, -19, -18, -15, 25, -46, -61, 18, -1, -23, -16, -49, -15, -26, 13, -15, 12, -54, -61, 2, -8, 5, -35, -32, 27, -20, -19, -11, 7, -66, -82, 26, -6, -6, -29, -13, 5, -3, -37, 13, 18, -9, -64, 12, 10, 3, 3),
    (30, -23, -3, 0, -14, 20, 9, -1, -24, 5, -15, 14, 18, -22, -5, -2, -13, 22, 16, -2, -17, 4, 2, 2, 6, -14, -16, -1, -4, 14, 25, 6, -21, 6, -14, 4, -3, -9, 6, -17, -27, 14, 7, 1, -45, 3, 3, -13, -15, -10, 6, -6, -44, 7, 34, -10, -11, 10, -10, 10, -1, -17, -7, 6, -14, 16, 14, -6, 17, 16, 10, 4, -11, 3, 7, 17, -3, -6, -30, 2, 14, 0, 11, -7, 5, 2, 6, 14, -7, -16, -29, 13, 16, 5, 12, 7, 6, -5, 17, 4, -12, 10, -26, 5, 2, 15, 16, 7, -9),
    (-52, 4, 3, -22, -3, -16, 7, -14, -38, -8, -11, -34, -51, 13, 1, -27, 2, -5, 4, -6, -24, -6, -2, -45, -10, 10, 4, -16, 1, -12, 10, 1, -30, -10, -12, -25, -7, 9, 16, 20, -1, -4, 16, 5, 21, -11, -1, 22, -21, 17, 18, 11, 21, -17, 20, 3, 4, 8, 17, 17, 2, 7, 17, 13, 15, -6, 12, 2, -18, 6, 6, 17, -2, -12, 6, 8, 1, -7, 9, -2, 15, -12, -8, 4, -10, -13, 10, 10, 14, -18, 27, -6, 21, -14, -2, -4, 3, -2, -11, 3, 7, -2, 14, -5, 7, -10, -3, 6, -5),
    (1, 2, -4, 17, 3, 2, -3, 5, -19, -2, 2, 9, 2, -8, -14, 21, -7, -10, -18, 10, 1, -6, 3, 2, 4, -8, -16, 5, -14, -7, -10, -1, 7, 5, 13, -8, 6, 2, -23, 15, -2, -4, -6, 2, -15, -13, 5, 7, -2, 3, -14, 15, -3, -11, -23, 18, -29, -6, 12, 8, -7, -2, -9, 0, -1, -14, -17, 18, -12, -4, 12, 2, 9, -3, -6, 12, -8, -4, -2, 5, 2, 10, 13, -5, 10, -9, -10, 12, -3, -2, 2, 16, -10, -6, 2, 6, -2, -8, -2, 15, 0, 2, -6, 8, -10, 0, 16, -2, -3),
    (13, -9, -3, -3, -8, 16, 15, -7, 23, 3, 2, 1, 20, -17, 14, 1, -15, 19, 28, -3, 4, 25, 19, 11, 2, -14, 10, 13, 0, -1, 12, 0, -3, 15, -8, 6, 1, -14, 22, 7, -10, 1, 20, -6, 13, 7, 19, -2, 27, -27, 18, 7, -30, 23, 31, -3, 26, 23, 0, -7, 18, -16, 8, 3, -2, 17, 20, -2, 15, 19, 4, -2, 10, -6, 1, 13, -10, -2, 11, 2, 6, -9, 3, 11, -3, -8, 17, -11, -6, 13, 9, -2, -12, 14, -2, -3, -2, -4, 16, -1, 1, 2, 9, 6, 2, 3, -2, 0, 0),
    (2, -3, -4, 15, 2, -14, -6, -7, 9, 2, 13, -15, 5, 1, 6, 8, 6, -10, -7, -7, 7, 6, 3, 3, -2, 15, -13, 10, -3, -3, -8, -2, 2, -5, -6, -9, -14, 6, -20, 19, 26, -18, 7, -6, 13, -11, 9, 8, -9, 22, -11, 10, 27, -18, -23, 0, 11, -7, 5, 7, -17, 22, -14, -5, -1, -17, -12, 10, 7, -10, 19, -1, 2, 2, -10, 2, 4, -7, 6, -15, 10, -1, -19, 10, -3, 22, -13, 7, 12, -9, -7, -6, -2, -1, -3, 5, -2, 9, -2, 2, -16, 5, -3, -10, 7, 6, -3, 14, -4),
    (-15, 4, 22, 18, -2, -6, 2, 14, -59, -3, 6, 21, -6, 3, 18, 11, -2, -18, 0, 13, 3, -7, 3, 18, -6, -10, -3, 10, 17, 4, 13, 10, 9, -11, 24, 12, -6, -12, 19, 8, -15, -10, -1, 6, -74, -14, -8, 6, -16, -3, 38, -4, -5, -34, -15, 18, -14, -45, -17, 3, -5, -2, 18, 10, 20, -14, -7, 14, 17, -38, 3, -1, 16, -9, 15, 0, -24, 9, -6, 3, -28, -2, -21, -4, 5, 8, -7, 2, -6, 6, -7, 5, -18, -27, -34, -2, 0, 9, -22, 1, 13, -6, -5, 0, 9, -35, -38, 1, -1),
    (-27, -20, -11, -33, 8, -20, -24, -14, -53, -12, -14, 0, 10, 3, 7, -7, -6, -5, -29, 16, 40, -10, 3, 4, 18, 6, 15, 3, -16, 11, 14, 22, 5, 3, -1, 10, -34, -46, 8, -39, 1, -17, -32, -34, -33, -1, -18, -16, 22, -5, 6, 14, -23, 3, -46, 26, 33, -5, 2, -9, 10, 10, 21, 12, -15, 25, -2, 29, 18, -6, 14, -2, -12, -24, 2, -30, 2, -18, 0, -41, -8, -9, -1, -23, 11, 4, 9, 11, -14, 7, -8, 22, 20, -2, 10, -8, 8, 11, 4, -8, -5, 22, 7, 30, 11, 4, -6, 9, 0),
    (-17, 20, 1, 2, 12, 1, -18, -1, 11, -6, -15, 7, -12, 7, 19, -12, 9, 5, -8, 10, 9, 1, -3, 16, 7, -14, 14, 3, 19, -3, 10, -1, -6, 18, 5, 27, -26, 35, -14, -14, 31, -5, -21, -6, -35, -14, -8, -19, -26, 42, -18, -16, 35, -6, -32, -16, -34, -25, -25, -24, -6, -20, -20, -22, 23, 8, -25, -19, -6, -1, -6, -9, 24, 19, 5, 20, -7, 15, -6, 18, -19, 4, 11, 2, 4, 17, 7, 10, 4, -7, -13, 18, -44, -7, 8, 8, -5, -2, 0, 1, 2, -9, -24, 6, -22, -10, -5, -4, 0),
    (19, -9, 17, 2, -13, 17, 7, 8, -10, -1, -6, 18, 6, -11, 24, 14, -42, -6, -7, 6, 15, -15, -7, 1, -9, -26, -8, -15, -39, -33, 7, -21, 25, -74, -32, -7, 19, -3, 17, 22, -19, 26, 0, 25, -12, 9, 4, 19, 6, -3, 37, 8, -50, -4, -6, 21, -11, -11, -5, 6, 6, -5, -6, -14, -43, -24, 2, -9, 23, -42, -20, -17, 21, -6, 22, 17, -15, 36, -14, 28, 3, 9, -5, 2, 20, -6, 15, -1, -20, 5, 2, 23, -2, 10, 2, 4, 1, 3, -17, -16, -12, -10, -1, -14, 2, -2, -7, -21, 0)
  );
  ----------------
  CONSTANT Layer_4_Columns    : NATURAL := 16;
  CONSTANT Layer_4_Rows       : NATURAL := 16;
  CONSTANT Layer_4_Strides    : NATURAL := 2;
  CONSTANT Layer_4_Activation : Activation_T := relu;
  CONSTANT Layer_4_Padding    : Padding_T := same;
  CONSTANT Layer_4_Values     : NATURAL := 16;
  CONSTANT Layer_4_Filter_X   : NATURAL := 3;
  CONSTANT Layer_4_Filter_Y   : NATURAL := 3;
  CONSTANT Layer_4_Filters    : NATURAL := 24;
  CONSTANT Layer_4_Inputs     : NATURAL := 145;
  CONSTANT Layer_4_Out_Offset : INTEGER := 6;
  CONSTANT Layer_4_Offset     : INTEGER := 1;
  CONSTANT Layer_4 : CNN_Weights_T(0 to Layer_4_Filters-1, 0 to Layer_4_Inputs-1) :=
  (
    (1, -21, -2, 3, -13, -21, -17, -14, -12, -16, 2, -39, -17, 20, -21, 23, -10, -6, 5, 1, 10, -15, 14, 5, -4, -12, -3, -26, -19, 11, -26, 11, 11, -14, -4, 1, 10, -1, 9, -1, 9, 1, -2, 15, 2, -15, -8, -5, -13, -3, -2, -4, -5, -23, -25, -5, -16, -10, 1, -61, -11, 20, -17, 18, -6, -12, 2, 18, 10, 1, 7, 13, -15, 0, 6, -28, 23, 21, -23, 12, 18, -15, 0, 9, 12, -10, 22, 2, 8, 2, -2, 0, 8, -14, -8, 5, -1, -10, 15, 6, -1, -5, -2, 9, -2, 3, 18, -21, -1, 21, -14, 15, -4, -6, 12, 14, -9, 7, 11, 2, 3, -4, 18, -7, 21, 28, -16, 16, -1, -9, 3, 17, -3, 2, 26, 2, 10, -10, -7, -4, 6, -15, -6, -4, 1),
    (-6, 0, -6, -4, 15, -3, -6, 9, 7, -4, 0, 5, 0, 6, -7, -2, -2, 2, 6, 10, 19, 0, 3, 8, 8, 1, 13, -6, 1, 12, -10, -15, 7, -11, -5, 2, 6, -8, 17, -2, 9, -9, -16, 4, -3, 1, 3, -8, -31, 0, 15, 0, -10, 27, -26, 15, -6, 7, 14, -1, 2, 18, -56, -7, -22, 14, 7, 28, 6, 23, -30, 18, -12, 5, 11, 3, -2, 18, -42, -31, -12, 6, -11, 30, 7, -3, 3, 11, -1, -19, -2, 0, -17, -2, -2, -24, -9, 18, 3, -7, -3, 14, -29, -4, -19, 15, 2, 7, 0, 8, -13, 3, -13, 14, -1, -6, -6, 12, -38, 6, -14, 17, -6, 17, 3, 10, 4, -5, -2, -2, -10, 9, -2, 1, -17, 0, -2, 4, 5, 2, 2, -2, 10, -9, -11),
    (-2, 8, -2, -3, 3, 4, -3, -9, -2, 10, -3, 7, 7, -7, 13, -18, 25, 15, -7, -14, -4, 12, -7, -5, 4, 6, 2, 8, 14, -10, 3, -6, 24, 22, 3, -6, 1, 10, -3, 3, 10, 14, 18, 14, 17, -11, -2, 0, 18, -24, 6, -3, 19, -20, 18, -15, -3, -27, -9, -34, 3, 10, -8, -27, 10, -10, 19, 4, 27, -12, 11, -23, -13, -8, -13, -16, 3, 1, -6, 7, -1, -14, 21, 10, 22, -4, -2, -22, -18, -6, -13, -14, 5, 5, 0, 8, -18, -15, 7, 6, -4, -12, 14, -3, 4, -19, -14, -20, 21, 0, -10, -39, -17, -10, 4, 19, -26, -4, 2, -2, -3, -16, -3, -19, 9, 1, -1, 3, -4, -25, 7, 7, -15, 2, 13, -7, 6, -22, -7, -14, -9, 5, -11, 2, -2),
    (-6, -1, 2, -2, -6, -14, -7, 6, -6, -18, 2, -2, -1, 0, 6, -2, -7, -3, 20, -5, 16, 13, -10, -7, 7, 12, 24, 4, 6, 23, -17, 14, -36, -31, 0, -5, -9, -1, -12, -10, 4, -11, 6, -10, 1, -8, -13, 17, 1, 1, 8, 1, -11, 2, -9, 7, -7, -7, 11, -4, 9, 6, 0, 0, -7, -5, 23, 8, 4, 5, -22, -12, -15, -2, 14, -4, 11, 34, -10, 22, -28, -38, -48, -2, -18, 10, -41, -27, -30, -12, -15, -1, 9, -2, -13, 11, -2, -4, 10, -1, -6, 2, -3, 3, -1, 2, 2, 7, 0, -10, 0, -3, -6, -1, 10, 4, -10, 9, -24, 0, -5, -3, -6, 1, -8, 10, 1, 5, 4, -27, -33, 9, -10, 13, -8, -12, -3, -19, -26, 18, -7, 1, 10, -5, 6),
    (-6, 10, 1, -11, 5, -11, 11, -12, -5, -40, -15, -16, -15, -15, 8, 1, 13, 18, 4, -16, -6, -16, 17, -11, 4, -11, -1, 0, -11, -7, 16, 27, 11, 10, 16, -13, 3, 2, 7, 7, 6, 17, 12, 14, 1, 10, 10, 32, 3, 4, -11, -21, -35, -27, 10, -10, -12, -37, -18, -15, 12, 5, 25, -1, 21, 12, -11, -13, -15, -24, 39, -10, 11, -6, -5, -7, -15, -21, 30, 11, 15, 11, 12, -2, -2, -5, 26, 6, 22, -1, 11, 5, -11, -6, 12, 18, 6, 2, -7, -4, -32, -7, -6, -5, 1, -4, -10, -14, 23, 9, 9, -4, 19, -5, -15, -7, -24, -10, 22, -4, 6, -3, 2, -10, 8, -14, 23, -4, 11, -2, -3, 5, -2, -9, 13, 2, 15, 0, 11, 1, -2, -16, 12, -2, -4),
    (-4, -2, -6, -1, -3, -9, -10, 1, 6, -2, 6, 1, -2, 24, 9, 17, 12, 2, -28, 3, -13, -5, -4, 10, 6, 4, -2, -2, -2, -6, 15, -7, 11, 17, -12, -2, -11, -3, 7, 15, 9, 9, 8, 4, 10, -14, 3, -1, 8, 4, -27, -4, -11, -24, -14, -4, 2, -9, -25, -6, 4, 1, 12, 11, 26, 8, -23, -21, -10, -13, 0, 2, 18, 3, -14, 8, 10, -6, 26, 11, 15, 7, -11, -14, -7, -9, 8, -5, 27, 3, -1, 9, 18, -11, 11, 12, 11, 9, -14, -16, -5, -32, 3, -13, -6, -32, -25, -14, -14, -29, 12, -8, 6, 10, -2, -23, 6, -15, 12, -9, 14, 0, -10, -2, -22, -22, 20, 14, 3, 12, 2, -4, 15, -9, 10, 2, 16, 6, 8, 7, -11, 3, 12, 21, 1),
    (-12, 1, -8, -12, -43, -30, -35, -13, -12, -30, -14, -9, -5, 0, -6, -5, -3, 12, -22, -18, -26, 3, -42, 0, -29, -14, -18, 2, 6, 6, -2, -3, -25, 22, -8, -11, -12, 25, -21, 1, -10, 10, -2, 0, 14, 8, -3, -5, 15, 4, -9, -8, -5, 2, -20, 13, 5, -6, -11, 9, 29, 1, -4, -31, 14, 3, -27, -3, -15, 6, -27, 0, 2, -11, -23, 22, 11, -7, 13, -17, 9, 4, -21, 6, 1, 6, -3, -2, -2, -12, -16, 6, 0, -24, 13, -6, 10, 8, 2, 3, 9, 10, -22, 5, 10, 5, -2, 11, 0, -6, -3, -12, 18, 10, -3, 1, -2, 12, -9, 11, 21, 6, -10, 17, 8, 1, 15, -16, 18, -2, -2, 3, -6, 10, 16, 11, 23, 12, -7, 8, -2, -3, 20, -7, 9),
    (2, 12, 2, 0, -1, -2, 1, 1, 2, 9, 7, 4, -8, -10, -14, -6, -3, 13, -1, 0, 1, 8, 2, -1, -8, 4, 5, 10, -19, -7, -14, -1, -9, 14, -3, 8, -1, 7, 4, 6, 3, 14, 11, -5, -2, -2, -9, 2, 8, 14, 2, 6, 10, -6, 6, 10, 2, 5, 2, 10, -12, -14, -2, -10, -4, 7, -4, -2, 15, 2, 4, 9, -2, 11, 2, 10, -17, -18, -6, -6, -6, 10, 0, -2, 18, 6, -5, -4, -2, 5, 0, 12, -10, -14, -5, -6, -5, -4, 4, 3, 1, 6, 2, 4, 2, 11, -5, 2, -14, -1, -4, -6, -3, 6, 11, 4, 12, 8, 1, 11, 6, 10, 10, 9, -10, -8, -14, -14, 2, 3, 6, 6, 2, 4, -1, 0, 5, -2, -3, 9, -2, -1, -10, -6, -7),
    (8, -7, -2, -6, 2, -15, 13, 12, 14, 3, 6, -2, -18, -10, 10, -15, -6, -1, -7, -2, 22, -26, -5, 5, 5, -2, -2, -7, -36, -10, 16, 0, -12, -22, 3, 6, 22, -17, -9, 10, -10, -1, -6, -5, -37, 0, 26, 14, 11, 9, -10, -7, -2, 15, 9, 21, 21, 14, 13, 14, 19, 2, 6, -9, 21, 10, -17, 1, -15, -5, 6, 27, 16, 2, 13, 9, 22, -4, 0, -14, 11, 14, -6, 1, -15, -10, -14, 12, -4, 10, 14, 4, 6, 2, -6, -5, 5, -6, -5, -4, -3, 10, 1, 0, 6, 8, 5, 3, 18, 6, -6, -4, 20, -2, -13, -8, 2, 2, -2, 2, 21, 3, 0, 1, 32, 2, -5, -10, 18, -7, 0, -5, 4, -9, -5, 1, 15, -6, -6, -2, 17, -8, 3, -2, -2),
    (-9, -4, 9, 3, -2, 11, -3, -10, -3, 10, 4, 2, 6, -17, -15, -2, -22, 1, 4, -2, -3, 6, -11, 10, -10, 8, 0, 8, 10, -3, -18, -8, -3, 9, 2, -6, -2, 9, -14, 4, -4, 7, 10, -4, 11, 6, -15, -9, -7, 15, 6, -15, 4, 1, -12, -13, -17, 10, 10, 6, -7, -9, 6, 8, -17, 19, 6, -25, -9, 10, -31, -6, -18, 20, 12, 2, -4, -7, -24, 11, -8, 7, 2, -7, -5, 12, -22, 1, -10, 13, 9, 3, 6, 10, -22, 2, 8, 4, -1, -5, 9, -2, -11, -3, -2, -9, 2, -2, 5, -11, 10, -2, -4, 14, -1, -1, 2, 7, -11, -10, -9, 6, -6, -2, -11, -14, -1, -2, -9, 18, 2, -11, -1, 12, -3, -3, -12, 21, 4, 8, -1, -2, -10, -1, -5),
    (-14, 1, 14, 10, 15, 4, 14, 12, -14, -6, 13, -13, -3, 14, -11, 5, 12, 1, 22, 28, 22, 4, 5, 15, 8, 7, 22, 6, 7, 10, -24, -2, 10, 5, 12, 17, 7, 4, -12, 7, -3, 3, 6, 2, 11, -1, -23, -10, -19, -6, -11, 18, -8, -2, 9, 28, 6, -13, 6, -13, 20, 12, 3, -4, -22, -13, 3, 17, 17, -8, 9, 2, 14, 1, 9, -14, 6, 7, 0, -17, -7, -10, -4, -9, 13, -16, -5, -6, -7, -3, -1, -14, -5, -5, -3, -19, -43, -3, -11, -16, -18, -10, 8, -18, -7, -17, -25, -10, 21, 5, -14, -38, -27, -9, 10, 3, 9, -25, 12, -9, -18, -11, -3, -15, -6, -15, -17, -25, 7, -12, 10, 2, -9, -19, -9, 12, -11, -19, -3, -15, -5, -1, -21, -7, -5),
    (6, 6, -2, -18, 6, -6, 5, -6, 7, 4, 1, 8, -9, -9, -9, 5, 6, -2, 12, -7, -10, -11, -7, -8, 1, 4, 1, 6, -4, -16, -4, 10, -4, -2, 18, 11, -4, 6, 0, -2, 5, -1, 14, 3, 8, 4, -10, -5, -14, 4, 20, 5, 15, -6, 18, -5, 2, 11, 17, 1, -10, -6, -41, 9, -18, 1, 32, 7, 10, 2, -6, -14, 1, 14, 14, -1, 16, -2, -44, 10, -37, -15, 6, -12, 9, 11, -14, -24, -6, 14, 8, 9, 23, 5, -15, 6, -32, -1, -4, -10, 4, 1, -1, 5, -16, -7, 14, -6, 0, -5, -24, -6, -52, 4, -5, 0, 4, -10, -24, -6, -35, -17, 11, -3, 2, 0, -14, -4, -50, -7, -26, -8, 9, -7, -10, -11, -33, -6, 5, 5, -2, -2, -8, 6, -3),
    (1, 2, -2, -24, -19, 14, -8, -13, -7, -6, -19, 20, 7, 3, 26, 13, 4, -2, -13, -23, -22, 6, -50, -7, -15, -9, -23, -3, -21, -6, 6, -2, -4, 14, 23, 0, 7, 6, -14, 4, -3, 10, 18, -5, -2, 6, -13, 4, 6, 5, -6, -17, -28, -41, -10, -15, -10, -10, -27, -18, -19, -16, -2, -11, -42, -2, 23, -7, 7, 16, -40, 13, -12, 5, 15, -22, -7, -2, -40, 0, -38, 16, 16, 13, 10, 25, -26, 11, -11, 6, 11, 5, 17, 16, -31, -2, -40, 6, 9, -14, -27, -25, -13, -4, -15, -20, -7, -20, 15, -8, -22, -39, -48, 7, 9, -3, 6, 19, -43, 8, -35, 0, 3, -5, 7, 13, -24, 9, -23, 0, 3, -1, 0, 2, -22, 17, -13, 9, 6, 14, 8, 11, -5, 10, 1),
    (12, -9, 3, -11, -1, -9, -24, -15, -4, -4, -7, 3, -8, 2, 5, 8, 22, -4, -7, -10, 9, -21, -34, -4, 15, -2, -15, 4, 8, 5, 21, 10, 18, 5, -18, -8, 4, -9, -14, -16, 6, -12, -26, -8, 7, -7, 9, 3, 6, -3, 17, 6, 22, -10, 6, -8, 10, -5, 12, 0, -26, 4, -1, 21, 24, 0, 5, -7, 32, -6, 13, -4, 27, -2, -8, 6, -8, -24, 23, 12, 32, 9, -15, -28, 5, -10, 25, -1, 26, -4, -11, 13, 4, -29, 26, -1, -10, 0, -2, -15, 1, -2, 1, 6, -14, -21, 11, -2, -12, 16, 6, -1, -9, 6, -3, -5, -6, -2, -3, 11, -2, -17, 19, -7, -43, 10, 13, -7, -19, 5, -10, 4, 11, -7, -12, 15, 4, -10, 18, 3, -32, 2, -6, 2, -2),
    (3, -6, 17, -3, -1, -37, -6, 1, 0, -8, -31, -19, -17, 6, -3, -6, 15, -12, 22, 15, 16, -4, 18, 12, 13, -5, -6, -10, -8, -3, -17, -6, 16, -6, 12, 6, 10, -4, 14, 10, 10, 6, 4, 8, 7, -14, -10, -2, 14, -2, 26, 26, 14, 14, 17, 23, 18, 2, 27, -9, 10, 19, -11, -4, 14, -1, 18, 56, -2, 20, 4, 16, 13, -8, 0, 17, 29, 21, -12, -24, 6, -6, -5, 6, -4, 5, 1, -8, 10, -6, -17, 13, 6, -23, 10, -16, -10, 9, -3, 1, 2, 10, -16, -3, 7, -6, 2, 10, 1, 17, 17, -4, 3, -5, -34, -17, -12, -6, -4, -6, 6, -18, -23, 3, 6, -18, 32, -26, 9, -14, -38, -26, -10, -11, 1, -16, -1, -11, -38, -7, -13, -2, 14, -3, -1),
    (7, -9, 10, 3, -3, 18, -11, -3, -2, -6, -6, 9, 6, -5, 20, -13, -2, 0, -2, -14, -16, 22, -5, 5, 9, -2, -17, 5, 5, -29, 14, -12, 9, -2, -14, 11, -14, 9, 20, 17, 18, -2, -2, 8, 5, -65, 0, -6, 3, 7, 3, -20, 0, 2, 10, -9, -7, 4, -8, 6, -27, -11, 13, -3, 1, 1, -30, -63, 3, 6, -18, -23, -16, 19, -29, -1, -22, -7, 30, 6, -4, -45, -86, -64, -22, -3, -37, -42, -9, 9, -37, -13, 7, -1, 12, 17, 9, 10, 6, -20, 4, 0, 26, 3, 3, 23, 8, 4, -9, -9, 8, 11, -7, 0, 5, -31, 10, 1, 28, -20, -14, 26, 10, -8, -26, 2, 5, 22, -41, -19, -3, -49, 22, -5, 18, -35, -19, 10, 17, -11, 9, 25, -12, 22, -11),
    (5, 17, 2, 27, 3, 16, -6, 19, 15, 14, 21, 9, 28, 13, -16, -1, 10, 14, 0, 41, -5, 7, -10, 18, 9, 3, 4, 18, 17, 15, -3, -14, -1, 5, -9, -1, -2, 4, -9, 3, 4, 2, 3, 10, 2, -18, 1, -12, -20, 6, -25, -10, -11, 15, -26, -2, 5, -8, -10, 20, 21, 7, 17, -20, 13, -12, -68, 7, -22, -1, -22, -12, 19, -11, -26, 9, 25, -14, 27, -30, 8, -19, -57, -6, -4, -13, 6, -18, 14, -6, -27, 2, 1, -52, 13, -17, 4, -3, -1, -23, 1, -9, 9, -20, 9, 2, -2, -1, -6, -13, 10, 0, 11, -14, -24, -11, 1, -9, -5, -20, 13, 0, -25, -8, 6, -24, 4, 7, 6, -32, -62, -25, -28, -1, -15, -27, 2, 4, -36, -4, -5, -16, -6, 7, 3),
    (-1, -4, 26, 9, 15, -4, 15, 6, 7, 6, 21, -4, -9, 6, -20, 17, -26, -3, 32, 14, 20, 9, 9, 18, 1, -15, 12, 0, -12, 17, -7, 21, -13, -6, 6, 6, 18, 6, 14, -1, 4, -14, 2, -6, -11, 6, 9, -3, -46, -25, 14, 1, 2, 2, 5, 11, -4, -17, 3, -2, 6, 14, -10, -2, -17, -24, 8, 9, -5, -22, -3, 5, -38, -26, 1, -27, -22, 3, -11, 6, 9, -18, 7, 8, 10, -16, 14, 1, -2, -20, 2, -34, -36, -4, -21, 7, 5, -18, 1, 5, -8, -9, 19, -6, -41, -7, -13, -6, 3, 4, -3, -2, 6, -17, 9, 3, 2, -24, 10, 13, 4, -7, -5, -40, -26, -4, -29, -2, 1, 0, 19, 14, 7, -2, 8, 12, 3, 0, 21, -13, 7, 10, -26, 18, -1),
    (-6, -27, -6, 14, -55, -16, -82, -24, -17, -5, -25, -17, -26, 6, -7, -6, -7, -32, -6, 13, -43, -12, -91, -18, -16, -13, -12, -28, -26, -2, 1, -10, -7, 3, -6, -3, -10, -19, -81, 1, -11, -10, -3, -14, 12, -14, 12, -2, -3, 4, -1, 2, -16, 14, -34, -6, -14, 7, 4, 4, 7, 22, -8, 22, -10, -6, -4, 1, -19, 11, -68, -7, -36, 20, 13, -10, 1, 29, -8, 24, -18, -13, -13, 5, -3, -4, -50, 5, -23, 11, 16, -23, -2, 12, -2, 9, 2, 6, -2, -3, -1, 1, -8, -11, -10, 11, 6, -6, 6, 9, 0, 31, 3, 9, 2, -2, 6, 14, -5, -6, -11, 19, 10, 3, 20, 29, 3, 26, -3, -11, 1, 0, 10, 6, 10, 2, -4, 6, 1, -4, 10, 16, -3, 6, -1),
    (-30, 10, 4, -15, -24, 14, -26, 2, -20, -1, 4, 6, -9, 11, -13, 8, -15, 13, 2, -2, -9, 23, -11, 3, -11, 5, 7, 2, -11, 6, -15, -21, -3, 8, -11, -2, 6, 6, -2, 6, -3, 1, 0, -1, -17, -5, -1, -14, -7, 15, 6, -9, -6, 8, -16, -18, -23, 16, -7, 6, 10, 1, -5, 3, -8, 18, -7, -15, -9, 28, -23, -26, -18, 25, -9, 14, 23, 9, -5, -14, 2, 3, -8, -23, -8, 11, 9, -16, 2, 10, -2, 3, 16, -12, 1, -10, -14, 3, 8, 6, 11, -14, -2, -9, -10, 2, 0, 6, -9, -1, -6, -25, -9, 6, 18, 2, 15, 2, 3, -37, -14, 16, -3, 3, -3, 6, 0, 1, -5, 1, 3, -27, 18, 3, 6, -32, -2, 8, -5, -4, 1, 6, -1, 6, -5),
    (-22, -11, 1, -5, 12, 22, -22, -11, -18, 18, 10, -5, 7, 23, -12, 6, -27, -22, -30, 2, -11, 5, -23, -17, -13, -1, -10, -26, 6, -12, 2, 8, 16, 2, -35, -25, 2, 7, 18, -12, 23, -5, -22, 3, 13, -36, -15, -20, -24, -6, 6, 2, 7, 14, -17, -16, -14, 12, 9, 1, -5, 19, -7, 11, -22, -14, -29, -3, -1, 4, -32, -9, -34, 11, -4, -19, -11, 23, 10, 14, -6, -26, -15, -10, 17, -1, -25, -17, 9, -23, -12, -7, -7, -25, 5, 1, -5, 10, 3, 8, 7, 14, -12, -6, -15, -1, -1, 3, -13, 15, -5, 12, -5, 12, 1, 4, -4, 8, -22, 4, -9, -3, -6, -5, 2, 13, -7, 10, -4, -24, -10, -7, 13, -10, 14, -12, -1, -20, 1, 6, -28, 7, -2, 8, 2),
    (14, -6, -23, 2, -35, -34, -26, -6, 8, -4, -50, -13, 2, -29, 12, -66, 17, -2, -19, -10, -14, -14, -2, 6, 4, 1, -37, 7, 4, -35, 9, -31, 18, -14, -11, -2, -17, -10, 11, 3, -23, -6, -13, -2, -17, -12, 4, -6, 4, -3, 3, 3, -13, -4, -20, -2, 1, -2, -14, 8, 14, -8, -6, -85, 18, 2, 3, 8, -3, -1, 10, 5, 10, 17, -14, 5, 14, -17, -20, -41, 18, 3, 17, 10, -13, -1, 6, 6, 11, 25, -6, -4, 25, -11, -15, -13, -19, 7, 12, 10, 1, 0, 4, -7, -13, 1, -1, -9, 3, -1, -27, -16, 0, 2, 16, 17, 18, -1, 8, -8, 2, 6, 7, 6, 6, -8, -27, -12, 6, 6, 16, 10, 8, 1, 7, 5, 12, 8, 8, 7, 10, 0, -2, -2, 3),
    (-8, -29, 3, 10, 7, -10, -7, 1, -15, -3, 4, -52, -17, 2, -25, 5, -15, -37, -6, 13, -8, -32, -6, -1, 2, -30, 4, -58, -57, -6, -1, 11, 3, -25, 5, 2, -17, -19, -3, -5, -7, -7, -1, -27, -8, 6, -1, 7, 8, -4, -1, 11, 2, -8, -5, 10, -16, 1, 2, -18, -20, -4, -10, 2, -5, -10, 4, 16, 17, -11, -1, 6, -19, 2, 18, -34, -6, 3, -30, -2, -16, -18, 16, 6, 2, -14, 15, -7, -20, -3, 6, -25, 2, -2, -35, -2, 14, 10, 4, 14, 6, 19, 11, 14, 15, 10, 13, 6, 10, 6, -6, -10, 6, 5, 10, 23, 6, 19, 2, 16, 2, -2, 15, 0, -10, 9, -26, -19, -11, -1, 2, 18, 2, 1, -8, 4, -16, -2, 9, 8, -7, 9, -22, -15, 0),
    (-2, 6, 5, -12, 1, -12, -10, -3, -2, -2, 2, 7, 2, -7, -13, -4, -31, -4, 14, 5, 7, 18, -25, 1, -16, 12, 3, 1, 14, 15, -22, 18, -23, 6, 7, 10, 8, 15, -9, 1, -10, 16, 6, 4, 18, 14, -13, 20, -47, -4, 8, -15, 5, -18, -16, -18, -29, 8, 5, -1, 2, -2, -19, 26, -73, 2, -8, -2, -7, 10, -49, -10, -55, 14, -7, 11, 18, 19, -6, 22, -30, 0, 0, -3, -2, 1, -22, 6, -23, 6, -2, 9, 1, 26, 7, 7, -81, -1, -5, -15, -10, -6, -29, -8, -41, -15, -1, 7, -8, 2, -13, 2, -33, 5, -25, -28, -28, 6, -27, -6, -46, -3, -9, -2, -2, 6, 1, -10, -2, 11, -11, -6, -10, 7, -6, 9, -14, 8, -11, -5, 5, 2, -2, -10, 1)
  );
  ----------------
  CONSTANT Layer_5_Columns    : NATURAL := 8;
  CONSTANT Layer_5_Rows       : NATURAL := 8;
  CONSTANT Layer_5_Strides    : NATURAL := 2;
  CONSTANT Layer_5_Activation : Activation_T := relu;
  CONSTANT Layer_5_Padding    : Padding_T := same;
  CONSTANT Layer_5_Values     : NATURAL := 24;
  CONSTANT Layer_5_Filter_X   : NATURAL := 3;
  CONSTANT Layer_5_Filter_Y   : NATURAL := 3;
  CONSTANT Layer_5_Filters    : NATURAL := 32;
  CONSTANT Layer_5_Inputs     : NATURAL := 217;
  CONSTANT Layer_5_Out_Offset : INTEGER := 6;
  CONSTANT Layer_5_Offset     : INTEGER := 1;
  CONSTANT Layer_5 : CNN_Weights_T(0 to Layer_5_Filters-1, 0 to Layer_5_Inputs-1) :=
  (
    (-2, -40, -4, -15, 1, 12, 14, -17, -16, -27, -20, -22, -14, -11, -13, -15, -26, -17, -13, -3, 5, -9, 6, -10, -16, -30, 3, -13, 4, 11, 18, 3, 5, -26, 0, -11, -3, -14, 9, -2, -14, -1, 5, -11, 4, -19, -13, -8, -14, -20, -16, -6, 7, 13, 9, -3, -2, 3, 15, -17, -8, -5, -6, 8, -11, 8, 18, -4, -1, -19, -15, -10, 9, -1, 7, 20, 5, 6, 14, 2, 9, -7, 1, 19, 12, 17, 14, -3, -3, -7, -2, -11, -3, 11, 9, -14, 11, -5, 7, 12, 1, -8, 29, -13, 8, -3, 18, 30, 8, 9, 21, -8, 1, -6, -2, 1, 1, 23, 14, 9, 2, -2, 10, -4, 5, 3, 18, -8, 14, -4, 8, 14, -5, -2, 11, -2, 6, -7, 5, 11, 0, 15, 9, 8, 5, -7, -7, 6, 5, -8, 1, -17, -18, -7, 9, 6, 6, -5, 7, 9, 0, -1, 0, -12, -1, -6, -19, 9, 5, 0, -14, 5, 3, -6, -9, -15, -19, -9, 10, 6, 7, 16, 8, 9, 10, 6, -6, -22, 2, 5, -14, 14, 12, -3, -2, -4, 3, 3, 0, -3, -7, -2, 10, 3, 1, 23, 5, 2, -2, 1, -1, -14, 2, 7, -6, 10, -2),
    (-19, -2, 6, -2, -1, -10, 23, -4, 1, -4, 9, 12, -9, -11, -1, 15, -7, -2, 1, 8, 2, 20, -6, -2, -29, -12, 4, 1, -7, -7, 14, 1, -6, -4, -2, 20, -24, -23, -6, 11, -39, -14, 19, 18, 11, 18, 6, -2, 2, 5, 11, -2, -3, -1, -16, -9, -1, 2, -22, -7, -2, -5, -4, 1, -27, -26, 21, 15, 9, -15, 17, 22, -2, 15, -34, 12, 2, -3, -1, 10, -5, 3, 9, 6, 10, 14, -6, 17, -23, 6, 1, -15, 19, 10, -18, -3, -6, 1, -30, 14, -3, 2, 5, 7, -20, 4, 20, 13, 0, 16, -14, 20, -56, -9, 7, -15, 21, 19, -29, -11, -4, 4, 2, -7, -9, -2, -14, -3, -9, 10, -16, 5, -11, -2, -9, 11, -33, -24, 7, 2, 16, -23, -14, -2, -8, 0, -3, 6, 8, 1, 1, 10, 6, 8, 2, 8, -13, 6, -11, 0, -1, 6, 9, 1, 5, -8, 2, -1, 1, 10, 8, 1, 7, 10, -27, 7, 2, 6, -1, 2, -18, -5, 0, -14, -4, 8, 0, 2, 7, -15, 4, -10, 5, 12, 4, 10, -37, -28, -14, -2, -4, -3, -2, -7, 0, -13, 19, -15, 1, -7, -11, -5, 9, -32, 14, -14, -7),
    (-4, 0, -13, -2, 1, -2, -10, 0, 0, 2, -6, -6, -3, -5, -9, -6, -15, -12, 14, -5, 18, -10, 6, -6, 13, 4, -37, 0, -3, -5, -22, -6, 2, 1, -23, -10, -2, 3, -12, -18, -33, -11, 22, -21, 6, -22, 12, -2, 14, 12, -28, 7, -6, 1, -3, -13, -4, -15, -12, -10, -2, 10, -7, -5, -10, 10, 2, -23, -8, -10, 6, -1, -8, 8, 38, 10, 3, 10, -17, 14, 7, 19, -10, -2, -3, -12, -4, -17, 4, -36, 22, 18, 0, -2, 1, -14, -1, 13, 37, 5, -3, 7, -27, 6, 7, 19, -24, 0, -10, -28, -9, -42, 1, -26, 22, 25, -15, -13, 11, -4, 6, 10, -1, 3, -8, 4, -9, -7, 10, 4, -20, -8, -4, -13, -3, -20, 11, -3, 3, 8, -7, -12, 15, -5, 1, -2, 2, 4, 14, 6, -6, 6, 2, 12, -7, -9, 10, -14, 3, -4, -4, -8, 4, 13, -3, -6, -16, 2, -2, 5, 7, 6, 14, 5, 3, 3, 2, 14, -4, -6, 2, -16, 8, 0, 5, -6, -11, 11, 4, -6, 2, -2, -10, 10, 1, 1, 2, 1, -3, 10, 2, -4, 1, -2, -2, -12, 5, -3, -3, -3, -5, 5, 2, 1, -2, 1, -23),
    (-8, -9, -11, -31, -13, 2, 4, -43, -29, -33, -37, -41, -8, 8, -33, -19, 1, -5, -8, -31, -1, -10, -13, -28, -1, -13, 12, 11, 13, 3, 10, -24, -18, -8, -36, -4, -11, 36, -50, -18, -4, -11, 27, -14, -1, -2, 5, 11, -6, -11, -6, 17, -7, 11, 0, -11, -6, 11, -8, 3, 1, 24, -24, -4, -2, -11, 12, 1, 22, -11, 4, 9, 22, -5, -26, 10, -13, 4, -14, -31, -34, 2, -25, -8, 6, -7, -11, -19, -30, -2, 16, -9, 4, 6, 15, 2, 16, -4, -17, 12, -5, -9, -27, -26, -20, 0, -8, 9, -3, 13, 1, -15, -11, 6, 32, -28, 10, -9, 19, 0, 7, -14, -9, 9, -5, -2, -7, -9, -14, 8, -6, -1, 10, 10, -6, -14, -3, -1, 18, 0, 6, -12, -10, 14, 19, -4, 3, 16, 5, 9, -7, 9, 7, 2, -14, 11, -1, -10, 9, -8, -8, 9, 19, 5, 6, -3, 22, -8, 18, 2, 3, -2, 4, -1, -26, 9, 2, 4, -16, -3, -2, -8, 8, -15, 0, 20, 17, 1, 5, -6, 26, -5, 5, 7, -10, -4, -1, -7, -14, 5, -4, 5, -20, 1, 6, -2, -4, 2, 0, 3, 3, -5, -3, -15, 10, 10, -1),
    (6, 1, 6, 2, 5, 10, 2, 7, 14, -5, -6, -7, -3, 6, 3, 14, 20, -10, -11, -2, 2, -25, 8, -5, -3, -21, -5, 20, -7, -21, 2, 11, -8, -7, 7, 14, -2, 3, -19, 4, -13, -3, -3, -2, 22, -17, -26, -37, -4, -27, -22, 4, -6, -9, -6, -28, -23, -13, -29, -5, -7, 10, -12, -3, -21, 12, 9, -26, 12, -4, 2, -37, 2, -8, 11, -8, -2, 14, 19, 1, 14, -11, 2, -24, -22, -4, 7, 11, 11, -15, -8, -2, -17, -28, 0, -12, -5, -18, 2, 0, 8, -13, -16, 5, -2, -17, 11, 9, -3, 1, 5, 12, -7, 14, -2, -23, 10, -14, -3, -49, 10, -15, -12, 11, 2, -15, -8, 7, -15, -17, 6, 4, 13, -4, 13, -8, 3, 14, -14, -29, 12, 5, 9, -31, -34, -17, 16, 1, 18, -2, 1, -11, -15, -15, -13, -16, -37, -23, -24, 12, -1, -4, -5, 1, -1, -2, -7, 17, 20, -18, -16, 5, -2, -11, -3, -4, -11, -10, -3, -3, 16, -6, -11, 10, -7, 26, -16, -13, 15, 14, 3, -5, 11, 10, -4, 12, -3, -10, -3, -2, 1, -9, -15, 6, 14, 3, 15, 2, 24, 11, -9, -2, 9, 3, 1, 24, 15),
    (8, -2, -27, 4, 8, 2, -18, 10, -6, -6, 2, -11, 12, 9, -10, 1, -13, 0, -6, -21, 8, -18, -14, 8, 6, -3, -30, 1, 5, 6, -15, 2, -10, -14, 10, -3, 10, 13, -1, 5, -11, 1, -13, -38, 11, -11, -18, -2, 7, 1, -37, 1, 3, 13, -7, 6, -2, 0, -7, 5, 14, 7, 2, 5, -6, 2, -8, -14, 10, 0, -7, 3, 6, 10, 15, -13, 4, -6, -35, 4, 14, 13, 12, 18, 2, -16, 2, -7, 18, -16, 9, 18, -10, -18, 9, 9, 18, 18, 16, -14, -8, -1, -21, 8, 31, 12, 14, 3, 2, -15, 10, -6, 21, -31, -9, 18, -15, -5, 16, 13, 1, 13, 1, -8, -2, 2, 11, 4, 14, 13, 6, -1, 2, -1, 8, -1, 6, -9, -39, 6, -1, 5, 11, 2, 1, -34, 5, -6, -1, -2, -16, -30, -36, -16, 17, -12, -9, -10, -5, 7, -7, 5, 18, -34, -27, -12, 6, -2, -33, -31, 9, -27, -23, -6, -24, -29, -29, -16, 11, -11, -18, -15, 2, 7, -5, 9, -10, -27, -17, -27, -15, 0, -41, -17, 2, -18, -42, -8, -8, -14, -57, -20, 2, -23, -33, 4, -21, 9, 3, 1, -30, -11, -15, -31, -19, -9, 10),
    (-7, -18, 9, -27, 6, 17, 3, -12, 6, -18, -16, -49, -18, 1, -1, -16, -22, -9, -5, -15, -67, -6, 14, -12, -28, -26, -18, -10, 12, 0, 4, 10, -2, 20, -25, -22, -11, -2, -30, -14, -7, -17, 4, 11, -50, -3, 2, -27, -4, 2, 4, 10, 2, -8, -16, 5, -12, 22, -5, 3, 5, -10, -14, -2, 4, -4, -13, 18, 13, -1, -13, -10, -10, 10, 12, -1, -10, -7, 12, -12, 13, 3, -14, -1, 3, 2, -11, 17, -7, -12, 0, 10, -36, 10, -6, 18, -8, 9, 1, -13, -5, 14, 16, 0, 15, -2, -17, -7, -5, 7, -9, 10, 11, -10, 6, 16, -32, 2, 0, 6, 10, -12, -27, 2, 10, 10, 9, 1, 4, -4, -3, 1, -9, -10, -2, -7, 7, 9, 13, -2, -5, -22, 9, -24, 4, 0, -11, -2, -7, -13, -3, 2, -5, 7, 5, 14, 9, -1, -7, 3, -3, 2, 6, 6, 5, 14, -2, 14, -4, -2, 5, -8, -20, -14, 10, -7, -9, 4, 2, 13, 4, 2, -6, 7, -7, -5, 15, 15, -9, 17, -15, 19, -13, 2, 16, -15, -19, 5, -22, -17, 6, -5, 9, -1, -14, 0, 8, 10, 1, -7, 6, 9, -4, -10, -27, 7, -7),
    (6, -7, 5, 11, -3, 3, 15, -9, 0, -1, 3, 6, 0, 6, 14, -3, -7, 2, 5, -23, 5, 4, 19, 6, 12, -13, 8, 13, -6, 10, 13, -9, -5, -7, 8, 6, -6, 18, 11, -2, -30, 12, 8, -16, 12, 1, 5, 1, -5, -1, -1, 6, -4, 10, 9, 1, -6, -3, -10, -6, -4, 14, -2, -1, -14, 0, 3, -2, 8, -10, -10, -8, 7, 7, 1, 1, -9, -1, -2, 6, 13, -4, 3, -6, 6, 14, 6, -11, -1, 11, 2, -12, -8, 6, 6, -4, 18, 22, -9, 4, 0, -15, -35, 11, 0, -7, 6, -6, 13, 11, 2, -35, -11, 22, -12, -8, 2, -6, 6, 10, 16, 16, -4, 6, 2, -4, -23, 11, -6, 5, -5, -3, 22, -2, 6, -19, 5, 10, -28, -10, 1, -7, 6, 7, 8, 16, -6, -6, -10, -7, -6, 9, 6, 6, 0, -2, 16, -3, 10, -11, 8, 1, 3, 7, -6, -9, 13, 3, 14, 9, 17, -14, -6, -17, -4, 6, -2, -1, -1, -15, 30, -5, 6, -11, 22, -1, -10, 12, -20, -22, 15, 17, 6, -14, 8, -28, -8, -3, 6, -14, 0, -18, -6, -16, 13, -2, 6, 9, 16, -4, -12, 1, -11, 3, 0, 11, -15),
    (7, 4, 5, 15, 5, 10, 6, 18, -6, -2, 5, 9, 7, 13, -6, -11, -7, 17, -2, -16, 6, 0, 5, -12, 13, -2, 3, 18, 9, -3, -21, 6, -17, 2, 14, 22, 9, 4, 7, -30, -10, 29, 7, -28, 11, 27, 3, 15, -4, 12, -7, 22, -16, -8, 14, -14, -14, 2, 9, 0, -5, -6, 14, -18, 14, 23, 5, -12, 13, 18, -8, 7, 2, 11, 2, 7, 2, 14, -2, -6, -7, 3, 10, 4, 7, 24, 6, -11, 2, 13, -22, -16, 1, -26, 12, -9, -8, 8, -14, 25, -2, -7, 1, -12, -28, 0, -4, 9, 8, 6, -11, -23, -2, 7, -12, -13, 10, -7, -6, 21, 19, 13, -15, 8, 2, -5, 7, -17, -32, -14, -17, -10, 10, 4, 1, -16, -1, 2, -9, -10, 15, 20, -5, 2, -11, -16, -15, -1, -5, -4, -12, -13, -16, -8, -2, -9, -6, -6, -6, -8, -5, -1, -10, -18, -13, -56, -13, 7, -6, -8, -21, 7, -12, -20, -12, -14, -33, -16, -9, -2, 11, 3, -26, -14, -4, -1, -34, -7, 11, -30, -13, 6, -2, -11, -2, -6, 20, -9, -19, -20, -32, -25, 2, -7, 2, -16, 4, -12, -12, 6, -30, -23, 12, 12, -39, -12, 5),
    (19, 18, -15, -2, -75, -7, -41, -10, 3, -3, -17, -2, 19, -1, 13, -5, 28, 4, -8, 10, 5, -17, 13, 13, -28, -11, -14, 4, -6, -7, -5, -27, -6, -29, -14, -8, -1, 0, 12, 0, 14, -3, -16, -42, -5, 7, -6, -8, 0, -11, -8, 4, 9, -3, 2, -5, -14, 15, -7, 16, 8, -15, 8, -1, 6, 3, -1, 10, 1, 13, 0, 14, 6, -2, -10, 3, -1, -24, -18, 3, 9, 6, 1, 4, -9, -18, 8, 9, 11, -6, -5, 0, 18, -30, -3, -25, 11, -40, -1, -13, 6, 1, 7, -13, 1, -10, -10, 4, 7, -17, 6, 27, 4, 15, 1, 3, 11, 19, 5, 2, 11, 1, -8, 12, 2, -5, -14, -5, -8, 2, 7, 10, 21, -13, 13, 11, 20, 2, 3, 10, 19, 16, 6, 18, 7, 3, 4, -5, 4, -8, 0, 6, -6, 1, 9, 6, 7, -4, 17, 2, -4, 2, -5, 0, 1, 19, -5, -19, 7, 2, -10, 10, 0, -12, -8, -11, -2, 5, -7, 7, 13, -2, 15, -3, 18, -3, 2, 7, 9, 6, -2, 7, -15, 6, -3, 0, 2, -5, -2, -6, -3, -4, -9, -11, -13, -15, 11, 5, 20, -21, -8, 1, -2, -23, -14, -1, 5),
    (-2, -8, -5, -5, -3, -15, 8, 4, -2, -3, -2, 11, -12, -1, -5, 15, -4, -4, 11, -8, -1, 6, -1, -8, -7, -15, 4, 0, -3, -10, 2, -2, -10, 2, 2, 9, -30, -5, -5, 24, -8, -8, 13, -14, 9, -1, 13, -18, -3, -9, 1, 2, -19, -10, 0, -11, -14, -1, 1, 8, -11, 1, -13, 15, -3, -14, 6, -9, 2, 0, 13, 1, -15, 2, 26, 3, 5, 8, 11, 0, 6, 2, 14, 16, -14, -7, -13, -3, -3, 8, 12, -3, -1, 11, 4, 3, -22, -9, 44, 13, 5, 24, 16, 5, 17, 3, 14, 23, -21, 0, -19, -12, -19, 1, 17, -4, 19, 12, 8, 0, -12, -4, 19, 15, 0, 8, 2, -1, 12, 10, 8, 12, -11, -3, -14, -16, -23, -6, 12, 1, 10, -3, 15, 3, -11, -26, 0, 7, -1, 10, 4, -19, -16, -16, -7, -15, -5, 24, -6, -6, -14, -6, -20, -20, -1, 7, -15, -10, -5, -4, 10, 17, 1, 15, 14, 9, -3, -8, 3, 2, 0, 22, -15, 2, -19, 3, -15, -20, 16, 15, -7, 0, -7, 1, 2, 14, 10, 4, 9, 5, 2, -3, -6, 11, -3, 8, -14, -6, -15, 5, 2, 0, 3, 3, -1, 10, -2),
    (-3, 7, 10, -1, -3, -4, -28, 2, 4, 8, 2, 4, -2, -14, 1, -1, 2, -11, 7, 10, 2, -2, -7, 3, -1, 14, 19, -2, 0, -6, -14, 2, 19, 15, 6, 11, 3, -20, 2, -8, 8, -19, -3, 14, -2, 14, 10, 11, 0, 14, 12, -7, 0, -3, 1, 1, 14, 7, 0, 2, 2, -18, -5, -2, -1, -11, -18, 6, -4, 9, 23, 7, 8, -17, 8, 6, 12, -8, -20, -10, -27, -7, 14, -8, 5, -18, -10, -18, -24, 6, -6, -23, -37, 17, -2, -6, -2, -16, 16, 1, 8, -22, -37, -14, -54, -3, 14, 5, 14, -29, -2, -21, -10, 6, -16, -13, -3, 12, -29, 2, -6, -10, 4, 6, -2, -15, -35, -6, -33, -2, 8, 3, 6, -30, 12, -15, 2, -4, -20, -7, -3, -4, -21, -1, -3, -12, -8, 20, 22, 1, 24, -20, 0, -25, -2, -15, 8, -15, -7, 15, -7, 10, -11, 1, -11, 5, -3, 12, 4, -22, -7, 1, 19, -12, 22, -34, 2, -21, 1, -11, -2, -23, -8, -3, 5, 1, -2, -5, 5, -14, 1, 10, -5, -27, -22, 0, -14, -7, 9, -42, -17, -31, -5, -8, -47, 0, -21, -1, 6, -6, 12, -18, 4, -52, 11, -1, -13),
    (0, -17, 20, -10, 20, 8, 7, -10, -1, -9, -4, -1, -1, -2, 13, 2, -19, 1, 2, -17, -17, 7, 14, 18, -26, -7, 11, -20, 10, 12, -16, 2, 1, 1, 14, -8, -26, 6, -25, -18, -42, -14, 5, -18, -35, 0, -8, -1, -16, 5, -1, -6, 13, 12, -1, 12, 6, 19, -18, -8, -10, 6, -32, -2, -15, -25, 3, -7, -6, -1, -9, -11, -13, 4, -7, -4, 19, 2, 18, -11, 10, -26, -16, -6, -14, 4, 7, 5, 18, 3, -6, -11, -6, -4, 12, -5, -23, -25, -12, -28, 10, 8, 3, 2, -1, 15, -13, -22, -14, 2, -15, -27, -31, -5, 0, -21, -7, -6, -10, -20, -9, 1, -18, 5, 17, 6, -2, 17, -10, 25, -15, -5, 5, -8, -19, 0, -3, -18, -4, 14, 4, -8, -18, -7, -14, -1, -7, 4, -7, 1, -1, -18, 9, -2, -2, 12, -9, 0, -15, 3, 3, 10, -10, -30, 6, -8, -9, 5, -12, -5, -7, -27, 3, 14, 15, -6, 2, 11, -18, -15, 1, 7, -6, -1, 16, 2, 6, -4, -19, 0, -6, 0, 4, -7, -15, 19, 12, 5, -7, 14, -6, 11, -3, -4, 11, -7, -2, 2, 6, -14, 5, 2, -2, 1, -16, -8, 0),
    (1, 19, -10, -7, -2, -7, -2, 9, 6, 2, -6, -6, -7, 5, -2, 6, -18, 6, -16, -5, -1, -6, 4, -2, -10, 12, -14, 0, 3, -15, 4, 16, 6, -6, -6, -4, -10, 14, -12, 14, -19, 10, -13, -12, 2, -6, -2, -14, -1, 5, -20, 3, -8, -11, 0, -2, -6, -2, -1, -10, 5, 9, 0, 17, 3, 3, -5, -11, 1, -8, 6, -5, -15, 6, 9, -6, -8, 3, -1, 18, 6, 18, 9, 7, -5, 15, -16, 10, -19, -14, -9, 10, -3, 5, -8, 14, -18, 10, 26, 1, -4, 6, 13, 18, 7, 20, 9, 17, -15, 19, -23, 12, -22, -15, -6, 12, 3, 14, -2, 7, -9, 5, 9, 4, 3, 13, 14, 9, 9, 9, 7, 9, -1, -5, -8, 3, -7, -6, -1, 9, 3, 9, -2, 3, 4, 9, -16, -1, -3, -4, -9, -4, 0, -8, -3, -6, 3, -2, -3, -13, -7, 7, -4, 1, 2, -30, 8, 4, -2, 8, -15, -2, -7, -10, -19, 13, -11, 0, 7, 5, 1, 11, -7, -7, -15, 10, -11, 1, 9, -21, -6, 5, 3, 3, -2, 1, -6, -22, -34, 0, -8, -5, 7, 10, 6, -3, 10, -1, -3, 0, -6, 0, 10, -17, -10, 0, -6),
    (-3, 3, -1, -5, -10, -2, -1, -3, 13, 1, -4, 2, 3, -2, 6, 1, 5, -9, -6, 13, -3, -2, -3, -10, 6, 7, 4, -6, -13, -11, -19, 12, 2, 9, -8, 3, 16, -7, -2, -11, -3, -6, -13, 16, 1, 4, -5, -2, 7, 6, 13, 4, -9, -8, -11, 13, -9, 7, -2, -1, 17, -22, -4, -8, 0, 3, -17, 13, -1, 7, -3, -2, -2, 19, -6, -2, 8, -22, -29, 10, 6, 3, -1, 11, 31, -12, 10, 1, 12, -1, -22, 13, -2, 9, -14, 2, 18, 7, -8, -1, 10, -32, -25, 10, -15, 4, -7, -1, 50, -26, 25, 10, 29, -19, -28, 12, -2, -16, -23, 15, 13, -12, -12, -18, -2, -12, 2, -4, -9, -2, -10, -16, 9, -2, 0, 30, 20, -10, -7, -6, -5, -18, 7, 13, -9, -21, -10, -8, 13, -5, -11, 12, -2, 2, 5, 8, -10, -1, -10, 9, 8, -5, -8, -6, 17, -49, -23, -2, -2, -34, 6, -8, 6, 3, -25, -4, 1, -18, -3, 10, -41, 7, -14, 30, -10, -14, -6, 4, 21, -42, -6, -29, -12, -30, 8, -2, 2, 4, 10, -21, -8, -28, 0, 8, -24, 14, -16, 11, -3, 5, 17, -2, 19, -1, -6, -22, -4),
    (-5, -13, -41, 14, -13, -17, 19, -31, -14, -14, -33, -9, 12, -10, -27, -11, -20, 2, -2, -11, -2, 15, -6, 0, 15, 5, -9, 10, 2, -15, 7, -5, 2, 2, -8, 13, 14, -2, 11, -5, 10, 9, 12, 10, 8, 10, 7, 31, 9, 1, -7, 4, -2, -10, 1, -6, 6, 7, 7, 5, 3, -11, 4, 7, 15, 7, 15, 2, -10, 13, 9, 21, 7, -11, -19, 10, -2, -4, 2, -24, -23, 2, -32, 3, 12, -10, -18, -11, -18, -2, 14, 15, 7, 5, -15, 14, 14, 3, -13, -6, -13, 3, 11, -18, -2, -5, -31, -5, 6, 4, 1, 20, 26, 10, 13, 13, -14, -4, 16, 32, -8, 2, -7, -5, -13, 12, 8, 2, 13, -2, -12, -14, -7, 1, 11, 11, 21, 2, 2, 3, -13, -7, 14, 0, 6, -2, -11, 8, 2, -5, 5, -12, -9, 9, -10, -5, 2, 0, -21, -7, -11, -7, 13, 11, -2, -29, -16, 4, -1, -4, -9, -12, 1, 9, 9, -3, 5, -3, -19, -25, -26, -2, -18, 8, 7, -13, 6, 5, -22, -26, 4, 0, 3, -15, -14, 5, -16, 1, 5, 1, 9, -2, 3, -2, -37, -1, -11, 10, 6, -11, 11, -7, -3, -13, -2, -15, -8),
    (5, 10, 6, -10, -2, 4, 3, 1, 6, 10, 6, -1, 9, 3, -2, 2, 6, -16, 3, 13, 2, -11, 21, 23, 14, 4, 0, -14, -6, 9, 4, 6, 19, 14, 11, 0, 2, -2, -2, 15, 6, -24, -11, 10, -18, -2, 16, 16, 0, 3, -1, 2, 6, 7, 15, 7, 6, 13, 7, 8, 1, 1, -8, 2, -8, -8, -41, 3, -5, -3, -11, -5, 5, -28, 8, -15, -13, 8, 14, -17, -31, -20, -17, -31, -23, -4, -43, 14, -2, -21, 22, 12, -32, 13, 16, -4, -14, 7, 2, -34, -32, 8, 7, -5, -7, -14, -11, -30, -28, -1, -14, 6, 6, -3, 3, 4, -19, 2, 3, -15, -3, 1, -10, -18, -31, -16, -18, -11, -18, -22, 3, -9, -33, 14, 10, 4, 2, 22, 22, -4, -14, 4, -7, -25, 0, -3, -14, -9, -17, -14, -8, -20, -34, -24, -44, -11, 14, 14, 1, -12, -51, 1, 12, -8, 1, 11, 22, 2, 1, -3, 2, -14, -10, -15, -10, -25, -33, 0, -23, 0, 9, 23, -16, -6, -24, -15, 6, -13, 3, -6, 13, 9, 8, 12, 3, 0, 8, -7, 7, -19, -10, -21, -19, -10, -8, 14, -10, -10, -7, 6, 11, -7, 0, -9, 10, -9, 0),
    (-9, -19, 0, 11, 2, -13, 15, -41, 1, -24, -27, -27, 6, -28, -6, 9, -13, -13, 6, 5, -18, 8, 0, 12, 2, -18, 13, 33, 12, 4, 11, -18, 8, -23, 9, 13, 15, 2, 10, -4, -5, 9, -4, -12, 11, 17, 2, -3, 0, -19, 3, 3, 13, 3, 7, -2, 5, -3, 16, 14, -6, 4, 11, 5, -5, -1, 6, -11, 2, 14, 1, 0, -7, -24, 5, 3, 5, 13, 17, -7, -14, -6, 19, 8, -2, 13, -2, 22, -18, -20, 5, -14, 10, 14, -19, -4, -12, -22, 11, -1, 12, 15, 13, -3, -3, -11, 14, -3, -18, 27, -11, 20, -30, -3, 14, -34, 13, 15, -19, 1, 0, -15, -3, 20, 15, 6, -3, 2, 0, -2, 10, 3, -3, 8, -10, 6, -33, 1, 14, -31, 16, 11, -11, -4, -5, -1, -4, 9, 6, 13, 3, 10, 6, -2, 8, -7, -5, 4, 0, 0, -2, -6, 1, -11, 5, 0, -8, -10, 0, 10, -10, 10, 3, 3, -8, 10, 8, -2, 3, -5, -8, 8, -5, -14, -10, 4, 14, 2, 13, -2, 13, -2, -2, 8, 4, 5, 6, -5, -6, -1, -4, 3, -3, 6, -2, -11, -2, -18, 2, -8, 2, 9, 0, -4, 4, 6, -1),
    (6, -2, 1, 2, 2, 7, 13, -11, 13, -10, -6, -4, 8, 0, 18, -1, 14, 13, -14, 4, -18, 4, 19, -3, 8, 6, 3, -2, 7, 9, 5, 6, 18, -23, 0, -7, -18, 11, 14, -2, 15, 12, -17, -9, -7, 8, 30, -42, -14, 4, -8, 12, 9, -4, 0, 3, 0, -24, 2, -3, -10, 12, 10, -4, 2, 14, 0, -14, 18, -2, 9, -31, -11, 9, -1, -12, 6, 1, -3, -10, -10, -10, -24, -33, 8, -5, 5, 23, 4, -37, -14, -14, 5, -10, -1, 7, -7, -6, 2, -12, 10, 6, 7, -10, 10, -15, -14, -28, -6, 4, 6, 33, 16, -23, -16, -15, 5, -24, -18, -4, -7, -26, -16, 10, 2, -13, -6, -3, 0, -12, 10, 2, -27, 5, -9, 23, 7, 10, -12, -24, 2, -16, -10, -34, -5, -16, 7, 21, 14, -4, 2, 3, 14, -7, 7, 7, -13, -16, -6, -9, -7, -6, -5, 1, 20, -9, 17, -6, -9, -27, 11, 13, 10, -3, 3, -5, 10, -13, 10, 5, -18, -7, 0, -7, -5, -1, 9, -5, 20, -11, 13, -17, -12, 2, -3, -6, -17, -15, 8, -4, -14, -7, 24, 0, 13, 5, -6, -8, 8, 1, 6, -3, 19, -3, -5, -26, 12),
    (8, 13, 4, -5, -10, -9, 13, 6, 4, -6, -25, -15, 16, 6, 14, 13, 11, 6, -31, -6, 3, 0, 0, 2, -22, -9, 1, -23, -2, -8, 31, 14, 13, -2, -11, -13, 18, 10, 17, 13, 15, 0, -13, 1, -15, 4, -7, -2, -46, -22, -5, 7, -2, -27, 14, 4, 13, -10, 1, 6, -19, 0, -14, 5, 0, -6, 11, 5, -7, 8, -6, -26, 12, 27, -27, -8, -16, -13, -1, -2, 14, 2, -26, -24, 38, 12, -2, 3, -1, 0, -30, 7, -3, -5, -10, 8, -5, 13, -10, -23, -35, -15, 23, -2, 6, -23, -16, -22, 15, 23, 3, 14, 10, 16, -30, -5, -21, -3, -13, -22, -34, -26, 0, 5, -16, -10, 16, 2, 10, -14, 16, -10, -21, 19, 0, 10, 1, -4, -6, -21, 5, -3, -28, -29, 7, 8, -16, -4, 2, 3, 2, 8, -2, 15, 3, -2, 17, 8, -6, 6, -6, 1, -8, 6, -1, -2, -5, 1, 17, 8, -2, -6, -10, -6, 2, 5, 1, 3, -5, -5, 1, 7, 5, 9, 1, 4, -7, 4, 2, -1, -12, -10, -15, -6, 8, 1, -6, -2, -3, 0, 9, -4, 0, -5, -26, 3, -7, 7, -3, -10, 6, -8, -2, 4, -12, -6, -2),
    (10, -30, -65, 2, -1, -22, -25, -30, -21, -19, -18, -1, 3, -20, 8, -50, -17, 1, 4, -16, 1, 6, 5, -3, 9, -5, -51, 2, -14, -26, -20, -12, -19, -23, -8, -5, 9, -14, 3, -43, 10, 10, -7, -27, 0, 6, 14, 2, -4, -11, -24, 5, -14, -30, 6, -11, -10, -24, -1, -6, 16, -6, 3, -10, 9, 10, 1, 2, -10, 9, 10, 3, 16, 15, -21, -15, -7, -23, 1, 7, 8, -3, -23, -12, 19, 4, 24, -31, 14, 16, -8, 1, -3, -2, 17, 23, 16, 18, -26, -19, -26, -31, -2, 0, 10, 6, -25, -25, 26, 4, 25, 3, 13, 13, -16, -3, -26, -4, 19, 27, 12, 10, -23, -17, -16, -13, -2, -3, 8, 13, -19, -1, 21, 2, 14, 14, 19, 7, -3, -10, -22, 3, 9, 5, 10, 11, 2, -7, -8, 1, -4, -6, 7, 6, -18, -9, 3, 2, -9, 3, -3, -19, 7, 10, -8, -12, 0, 13, 12, 3, 7, -3, -2, 11, -9, -2, 11, 3, -9, 2, 5, 1, -10, 5, -2, -14, 3, 4, -21, -13, 4, 13, 5, 4, 7, -9, 4, 6, 0, 1, -5, -3, 4, 9, 0, -2, -3, -9, 2, -4, -5, 3, -7, 4, 2, 3, -3),
    (-25, -12, -13, -19, -8, 7, 20, -32, -9, -9, -46, -37, -14, 10, -14, -33, -39, -25, -18, 2, 3, -17, -22, 15, -1, 0, -2, 10, -26, 11, 2, 1, -2, 13, -40, -10, 9, -3, -10, -19, -26, 4, -19, 24, -11, -20, -1, 6, -2, 1, -9, 9, -18, -3, 13, 0, 5, -10, -3, -7, -2, 17, -6, 0, -30, -16, -6, 17, -1, -3, -16, 1, -4, -27, -1, 19, 7, -8, -6, -17, -18, -8, -17, -2, 1, -3, 8, 8, -33, 7, 4, -19, 2, 9, 10, -5, 14, 17, -24, 2, -9, -21, -16, 13, -21, 16, -2, 11, 39, -1, 11, -4, 6, 11, -25, 21, 21, 6, 0, 11, 1, 9, -9, -7, -7, -10, 6, 6, -7, -8, 4, 1, 6, 7, 5, 0, -6, -2, -13, 12, -10, 7, -13, -5, 3, 6, -13, 6, -12, -13, 2, -1, 6, -7, -9, -9, 16, 6, 18, -3, 17, 6, -20, -13, 8, 1, -1, 13, 8, 21, -1, -15, -12, -9, -1, 11, 3, 8, -11, -18, 35, 5, 15, 1, 14, -13, -17, -1, -9, -7, 5, 11, 2, 6, -2, -10, -3, -1, -2, 5, 3, 2, 2, -4, -5, 5, 10, 6, 2, -9, -2, 1, -6, 0, -1, 2, 0),
    (9, -5, 0, 5, 2, 4, -13, -6, -23, 2, 9, -7, 4, -1, -3, 11, -3, 9, 10, -10, 10, -9, -10, -5, 8, -14, 14, 4, -6, 4, -18, -3, -19, -10, 9, 3, -7, 9, 7, 17, 14, 2, 21, -10, 10, -6, 2, -6, 9, -13, 3, 7, -13, 1, -12, 1, -4, -15, -4, 11, 5, 5, 10, -6, 15, 3, 17, -3, 18, 8, 8, -3, -1, 12, -11, 2, 3, -10, -17, 9, 6, 0, -9, 0, -10, -12, -11, -2, -31, -2, 2, -10, -2, -22, 7, -7, 6, 9, -12, -15, -5, -8, -26, 8, -2, -3, -18, -2, -7, 2, -11, -3, -10, -2, 14, -18, -6, -28, 21, 0, 8, 11, -20, -6, -18, -16, -22, -2, -16, -6, -4, -7, -3, 11, -5, 11, -13, 1, 12, -17, -7, -9, 14, 4, -1, -1, 32, -11, -2, -1, -10, 18, 14, 15, 18, 11, -6, 3, 3, -14, 15, -12, 17, 2, -13, -3, 3, 11, 6, 11, 33, -14, -4, -1, -5, 11, 13, 19, 10, 8, -7, -3, 4, -30, 2, -21, 7, 8, -22, -13, 20, 6, -3, 6, 0, -10, 1, 2, -10, 14, 14, 6, -11, -3, -2, -8, -2, -19, 6, -5, -5, 6, -10, -10, 17, 2, -26),
    (-19, -14, 0, 12, 17, 7, -3, 10, -5, 10, 14, -6, -10, 0, -14, 8, -6, -14, -2, -7, 3, -12, -11, -13, -9, 7, 9, 14, 22, 6, -10, 6, 7, 19, -3, 0, 2, -1, -10, 23, -1, -19, -13, -4, 19, -6, -15, -2, 2, 5, 4, 9, 11, 3, -6, -2, 11, -6, -6, -3, -6, -1, -1, 11, -9, -4, 4, -1, 10, -2, 0, -3, -18, -5, 0, 16, 17, 15, -2, 7, 7, -4, 4, -17, -15, -2, 0, -5, 2, -6, -5, -5, -9, -17, -13, -28, -8, 1, -21, 26, 41, 9, -2, 13, 2, 10, 9, -9, -7, 1, 1, 7, -2, -6, -21, 0, 34, -20, -22, -34, -2, 6, -7, 5, 21, 6, -4, 1, 7, 6, 7, 1, -3, 10, -3, 11, -12, -5, -9, -2, 17, -7, -13, -10, -2, 11, 10, 1, 0, -4, 9, 5, 6, -4, 7, -7, -2, -1, 5, -6, 6, -4, -5, 4, -3, 7, -13, -1, 0, 3, -9, 10, 13, 0, 0, 8, 9, 3, 8, -6, -9, 5, 3, -5, 1, -4, -4, 2, 14, -4, -4, -19, 1, -1, -17, -1, 12, 3, 3, 11, 6, 5, 5, -2, -4, 9, 0, 0, 0, 4, -8, -2, 12, -1, -3, -18, -1),
    (3, 3, -17, 7, -20, -12, -16, -12, -19, -3, -19, -12, 14, 4, -15, -8, -3, 11, -17, 5, 5, -13, -6, 24, -2, 28, -13, -15, -24, -11, -5, 5, -3, 4, -16, -7, 17, 23, -10, 4, -1, 18, -25, 0, -18, -8, 0, 23, -2, 11, -16, -5, -6, -6, -8, 7, 2, 4, -14, -2, 5, 17, -4, 5, 0, 5, -9, 0, -6, 2, -8, -5, 0, 3, -3, -17, -10, -6, -12, -6, -10, 18, -15, -1, 5, -13, 7, 5, 15, -17, 1, 7, -6, -13, 6, 12, -10, 21, 11, -10, -12, 10, -9, 16, 16, 18, -13, 1, 2, -21, -5, 5, -5, -29, -3, 23, -2, -2, -1, 0, -7, 4, 15, -5, 2, 18, -10, 14, 2, 12, -1, 7, -3, -15, -6, 1, -17, -17, -8, 12, 3, 7, -10, -12, 5, -9, 9, -8, 5, 9, -14, 4, 6, -8, 1, 9, 10, 8, 19, 0, 10, -10, -3, -19, 5, 7, 17, -13, 1, -4, 5, 4, 11, -2, -7, 2, -19, 0, 6, 6, 10, 7, 2, -9, -14, -1, -14, 4, 10, 0, 13, -6, -12, -12, 3, 2, -2, -10, 5, -10, -11, -9, 0, 6, 0, -5, 6, 6, 0, 4, -9, 0, -3, -5, -7, 2, -13),
    (-27, -28, 11, 23, 0, 1, 9, -34, -44, -15, -17, -18, -5, -4, -50, 2, -1, -30, 5, -4, -3, 2, -23, -5, -7, -3, 6, 4, -11, 4, 18, -6, -11, -8, -5, -3, 2, 14, -33, 19, 18, -17, 9, 5, 5, -6, -9, 2, 10, 15, 7, -11, -10, 2, -1, 1, 6, -3, 2, -7, -2, 6, -12, 9, 13, 8, 10, 6, -14, -12, -1, -4, 1, -28, -33, 3, 3, 12, 8, -17, -22, -3, -44, -22, 9, -5, -42, 16, -38, -10, 5, -15, 7, -6, -29, -3, 4, -22, -5, 19, 1, -2, 8, -18, -13, 11, -48, -9, 11, 7, -46, -7, -2, -16, 18, 3, 11, -16, -29, 10, 8, 7, -2, 2, -6, 13, 3, -14, 10, -1, -14, 1, -4, 3, -32, -10, 3, -1, 23, 11, -8, -20, -6, 18, -2, -21, -19, 7, 6, 25, 9, -14, -15, 5, -1, -14, 14, -19, -16, 3, 8, 2, 6, -5, -5, -2, -17, -6, 5, -7, -2, 29, 15, 6, -2, -11, -10, 6, -6, 6, 9, -3, -18, -7, 9, -9, 32, 2, 21, -9, -10, 2, -2, 2, 3, 10, 10, 6, 8, -14, 1, 10, -1, 1, -3, 6, -18, -10, 8, 1, 26, 1, 11, -6, -3, -1, 3),
    (-8, 21, -11, -3, -18, -2, -1, 2, 6, -2, -18, -5, 6, 0, 2, 6, 6, 8, -13, 6, -10, -4, -11, 13, -8, 10, 6, -19, -20, 5, 1, -10, 12, -13, -5, -13, 13, 14, 2, -5, 27, 9, -17, -11, -24, 6, 7, 3, -11, -13, -8, -22, 1, 20, 7, 5, -8, -7, -3, -12, -9, 16, -4, -6, 2, 2, -3, -19, -21, -16, 14, -3, -21, -20, 0, 10, 22, -6, -1, 6, -15, 14, 13, 13, -7, -11, -14, 22, -3, -14, 19, 6, 22, -3, -7, 2, -19, 3, 14, 3, -3, 6, -17, 1, -13, 9, -13, 6, -3, -13, -34, 21, -22, -21, 18, 18, 13, -8, -4, 7, -26, 22, 8, -7, -22, -24, -23, -14, 2, -4, -44, -18, -24, -2, -6, 20, 0, -18, 2, 10, 2, -16, -7, 9, -4, -9, 11, 7, 3, 18, 6, -12, -1, 2, -3, -5, -1, 2, 9, 7, 10, -9, 10, 1, 4, 4, -4, -4, -21, -22, -3, 3, 19, 26, -1, 2, -8, 11, 1, 0, -20, 16, -12, 16, -9, -10, 10, 18, 14, 5, 4, -3, -29, -22, -12, -11, 2, 18, 1, 2, -1, -8, 9, -4, -16, 21, -23, 6, -9, -14, -3, -14, -2, 7, -6, -22, 0),
    (-13, -22, -2, -7, -13, -13, 13, 8, -21, 16, 3, 11, -24, 0, -11, 5, 1, -19, 12, 13, 12, -12, -4, -2, -4, -9, 17, -16, -31, 7, 3, -24, -16, -13, -6, -38, -17, -10, -10, 13, -11, -25, 0, 38, -10, -38, -4, 14, -9, -5, 6, -18, -23, -8, -39, -32, -15, -37, 13, -35, 15, 3, -6, -4, -1, -30, -15, -21, -10, -24, -8, -9, -1, -11, 13, 3, -11, 0, 19, -19, -10, 2, -3, 11, -5, -26, 13, 5, 3, 1, 10, 22, 5, 19, 6, 14, -2, -14, 0, 9, -1, 11, 16, -14, -8, 10, -35, 7, -11, -40, 7, 6, -6, -9, 14, 36, 12, 6, 8, 28, 6, 6, 11, 16, -22, -15, 2, -30, -15, -7, 19, -13, -14, -16, -17, 10, 8, -27, 0, 20, 7, -39, 3, -15, -6, 2, -24, 15, 1, 4, 5, 3, -10, 7, 1, 3, 2, 8, -2, 4, -14, -9, -6, -6, 7, 19, -9, 3, -10, -5, -2, 17, 6, 16, 8, 9, -11, 8, -3, 13, -1, 10, -12, 14, -38, -26, 13, -11, 21, 13, -14, 4, -7, -6, -3, 3, 2, 11, -7, 2, -10, -2, -15, 7, -39, 2, -7, 18, -32, -25, 14, 6, 23, 8, 2, 6, 10),
    (2, -1, 2, 10, 9, -5, -6, 6, 2, 10, -12, 9, -4, -10, 3, -14, 6, 1, 15, 2, 9, 3, -5, 14, -6, -4, -4, 11, 7, -3, 1, -19, -1, 1, -2, -3, -6, -6, 0, -19, 18, 6, 13, 9, 6, -5, -3, 28, -15, 1, -5, -40, -50, -2, -17, -27, 1, -28, -7, -31, -22, -13, 7, 5, 5, -32, -7, 9, -11, -25, 5, -36, -13, 11, -10, 10, 13, 10, 6, -10, -2, 10, -11, 2, -5, -4, -10, -19, 15, -7, 4, 10, 13, 0, -2, 26, 1, 5, 4, -6, 13, 0, -7, -29, -9, 2, -13, -25, 8, -9, 7, -17, 14, -6, 6, 14, 13, 13, 15, 42, 0, -32, -12, -13, -28, -22, -22, -29, -16, -34, -24, -27, -6, -12, 9, 8, 6, -20, -5, -1, -4, -13, 14, -15, 6, 5, -2, -10, -3, -6, 11, -3, -1, -3, -14, -12, 8, 8, 14, -14, 18, -7, -17, 7, 9, -7, 11, -1, 18, 4, 9, -10, 1, -12, 7, -8, 1, -16, -19, -22, 14, 6, 22, -28, 16, 4, -15, 1, 3, -2, 17, 9, 5, -2, -6, 1, -4, -13, 5, 9, -5, -13, 4, -19, 14, 15, 11, -36, -10, 19, -5, -34, 10, -8, 12, 13, -1),
    (16, -2, -2, -16, 2, -3, 3, 7, 1, -9, 8, 8, 10, 11, 10, 10, -7, 6, 2, -10, -23, 13, 2, -18, 9, 6, 10, -14, -7, -6, 13, 0, 13, 1, 6, 7, -7, 11, 10, 0, 2, 2, -7, -6, -23, 25, 5, -15, -5, 7, -2, 2, -8, -3, 8, 1, 15, 0, 2, 8, 3, 1, 7, 7, 9, -15, -6, -6, -9, 23, -3, -1, 8, 3, -25, 8, 5, -21, -16, -14, -23, 6, -5, 14, 10, -11, 2, -6, 6, 12, -14, -9, 2, 13, 1, 3, 13, 5, -10, 10, 0, -24, -21, -10, -20, 7, 9, 17, 12, -17, 4, -30, -2, 14, 12, -10, 6, 18, -5, 17, 6, -3, 4, 7, 9, -8, -15, -8, -18, 4, 23, 10, 6, -12, 2, -15, -11, 3, 15, -5, 1, 2, -13, 13, -10, 6, -9, 3, -4, 3, -20, 2, -18, 8, 2, 9, 5, -11, -11, -8, -3, -11, 0, -14, 6, -10, -6, 1, -7, 3, -2, 7, 0, 1, -21, -14, -22, 7, 0, 4, -5, -17, -9, -22, 5, -11, 2, -7, -5, -13, 2, 10, -11, -4, 4, 7, 7, -5, -3, -16, -23, -9, 5, 8, -8, -13, 2, -17, -1, 2, -4, -3, 9, -18, -18, 6, -3),
    (6, 5, 3, 22, 18, -6, -35, -11, -24, 6, 8, 2, 12, -22, 12, -14, -10, -2, -17, -14, 2, 26, 1, -2, 10, -2, -8, 3, 26, -19, -25, 2, -31, 14, 3, 15, 46, -44, 26, -6, 14, -12, -8, 6, 14, -3, -25, 15, -1, -19, 2, -3, -14, -8, -2, -10, -33, -1, -7, -10, -22, -19, 6, 7, 18, -9, -10, -9, -2, -24, -9, 1, -15, -46, 3, 3, 9, -1, 8, -15, -10, -27, -4, -17, -15, -30, -23, -26, 0, -12, -18, 3, -11, -5, -15, 7, -10, -19, 0, -26, 5, -7, 11, 2, 1, -25, 0, -10, -31, -26, -14, -10, 18, -7, -10, -3, -17, 6, 12, 5, -10, -24, 1, -11, -18, -23, 10, -3, -20, -33, 7, -7, -10, -4, -8, -17, 7, 5, -6, -14, -6, 6, 14, -28, 5, 14, 3, -7, -14, -17, -4, 4, 5, -9, -22, -10, 17, 11, 9, -2, 6, 19, -9, 7, -40, 9, 1, 5, 5, 14, 3, -16, -19, -20, 8, 0, 6, 2, -9, 4, 29, 2, 10, 6, 22, 7, -7, 7, -6, 14, 16, 14, 6, 6, -3, -21, -6, -6, 8, 6, 2, 2, -5, -1, 23, 2, 6, 10, 19, -3, -6, 7, -9, 2, 13, 16, -1),
    (-21, 10, 10, 4, -2, 22, 14, 7, 9, 7, -9, -9, -15, 2, -6, 11, -1, -42, -6, -1, 1, 1, 0, -2, -34, -4, 20, 9, 0, 30, 14, 9, 14, 6, -7, 11, -24, 8, -14, -9, -18, -28, -6, 2, 15, -1, -1, -2, -20, -7, 9, 7, 7, 18, -2, 5, 6, 10, -2, 10, -7, 11, -16, -18, -20, -10, -6, 3, 13, 4, -21, 3, -15, -15, 9, 20, 9, 11, -2, 5, -16, -8, -15, 6, -4, 0, 10, -22, -24, -4, -2, -15, 22, -6, 0, -5, 1, 4, 2, 22, 6, -10, -5, -8, -18, -12, -2, 11, 9, -2, 23, -43, -19, 36, -8, -27, 17, 17, -10, 11, 3, 4, -4, 15, 2, -36, -20, -11, -19, -12, 9, 9, 17, -26, 27, -16, 7, 30, -3, -21, 4, 17, -1, 3, 15, 6, -7, 2, 3, -10, -2, -15, -1, -1, 17, 7, 5, -15, 12, -20, 9, 3, 9, -11, 3, -5, 6, 11, 9, -7, -6, 7, -5, -18, -9, -15, -15, -2, 12, -7, 6, -24, 14, -14, 16, 1, 12, -9, -7, -18, 8, 6, -1, -6, -20, 5, -7, -26, 3, -15, -27, -20, -2, -1, -3, -23, -4, -3, 13, -12, 0, -10, -11, -13, -8, 2, -17)
  );
  ----------------
  CONSTANT Layer_6_Columns    : NATURAL := 4;
  CONSTANT Layer_6_Rows       : NATURAL := 4;
  CONSTANT Layer_6_Strides    : NATURAL := 2;
  CONSTANT Layer_6_Activation : Activation_T := relu;
  CONSTANT Layer_6_Padding    : Padding_T := same;
  CONSTANT Layer_6_Values     : NATURAL := 32;
  CONSTANT Layer_6_Filter_X   : NATURAL := 3;
  CONSTANT Layer_6_Filter_Y   : NATURAL := 3;
  CONSTANT Layer_6_Filters    : NATURAL := 32;
  CONSTANT Layer_6_Inputs     : NATURAL := 289;
  CONSTANT Layer_6_Out_Offset : INTEGER := 6;
  CONSTANT Layer_6_Offset     : INTEGER := 1;
  CONSTANT Layer_6 : CNN_Weights_T(0 to Layer_6_Filters-1, 0 to Layer_6_Inputs-1) :=
  (
    (-20, -2, -6, -31, -7, 11, -8, -14, -4, -2, -1, 12, -2, 12, 22, 13, 6, -10, -16, 9, -18, 14, -21, -7, 15, -4, -1, -6, 12, 11, 9, 0, -15, -23, -15, -1, -1, 5, 5, -37, 0, -10, 3, 18, -14, 4, 0, 1, -5, -15, 2, -2, 0, 8, -7, 0, -2, -12, -3, -10, -2, 0, 17, -1, -23, -21, -43, 9, 6, -8, 2, -27, 11, -15, -6, 12, -9, -17, 0, -21, 7, -19, -1, -4, -4, -20, -13, -4, -16, -18, -7, -2, 4, -3, 2, 7, 7, -11, -2, 9, -5, -7, -4, -4, -17, 4, 8, 24, 1, 9, -3, -2, -2, -6, -2, 3, 8, 6, 8, -12, 14, 10, -14, 12, 7, -6, 2, 19, 15, 2, 5, -2, -6, -14, 9, 9, 3, -7, 8, 19, 4, 10, 0, 7, -4, 6, -6, 2, 13, 10, -13, -14, 14, 13, -1, -9, 13, 21, 1, 20, 11, 2, -4, -18, -5, -4, 4, 12, 2, -19, 9, 4, 8, -6, -4, 1, 4, 6, -1, 4, 13, 7, -19, -17, -1, -8, -8, -17, 4, 13, -5, -2, -10, -4, 2, 0, -4, -10, 6, -12, 19, 4, -14, -3, 10, -7, 1, -5, -14, 1, 4, -10, -15, 1, -13, 0, -3, -18, -14, -16, -6, 0, -4, -2, -9, -12, -1, 5, 5, -22, 9, -13, 20, 11, -2, -6, 8, 2, -1, -1, -15, 6, 5, -11, -31, 20, -29, 5, 0, -13, -14, 6, 10, 1, 1, -5, -25, -4, -15, 5, -2, -23, -22, -17, 14, 2, -15, -12, -3, -2, -12, 6, -4, -4, -5, -9, -16, -3, -25, -20, -17, -15, -2, 8, 9, 1, -8, 5, 11),
    (-24, -3, -1, 10, -1, 0, -5, -10, 7, 4, -7, -7, 2, -18, 9, -4, -3, 5, -13, -14, -1, 1, 12, -15, -7, 3, -15, 7, 18, 5, 13, -20, -9, 2, 6, 19, -6, 3, -14, -8, 22, 5, -15, -11, -24, -26, 4, -8, -2, -3, -7, -31, 3, 1, 18, -2, -12, -5, -13, -15, 9, -1, 14, -11, 16, -14, -9, 30, 9, 4, -9, 0, 16, -1, -9, -6, -1, -27, 0, 12, 5, 2, -8, -28, 5, 7, 20, -1, -5, 6, -14, -3, 18, 13, 14, 2, 13, 6, 16, 1, -13, -2, 13, 0, 23, -19, 21, 7, 2, -2, -9, -4, 2, 3, -15, -15, -4, -6, 9, -3, -3, 8, 5, 6, 0, 4, 14, -4, 15, -18, 6, 19, -18, 2, -7, 7, 17, -4, 14, 11, -6, -10, -4, -21, -2, -2, -2, -13, 10, -24, 14, -11, -6, -9, 2, 4, 4, -6, 16, 1, 14, -7, -5, 15, -13, 8, -2, 10, 15, -7, 4, 0, 4, 2, -5, -5, 4, 0, -3, -14, 15, 9, 10, -4, -7, 14, -5, 5, -3, 2, 29, 7, 1, -2, -3, 11, -1, -15, 4, -18, 6, -11, 2, -4, 11, -5, -10, -5, -2, 9, -8, -14, -27, -4, -16, 0, -12, 3, -2, -4, 4, 9, 8, 7, 4, -6, 13, 10, -4, -15, -4, 8, 16, -5, 0, -3, 18, 6, -6, -9, -11, 14, -11, -16, -34, 5, -20, -2, -17, -5, 5, 12, 9, 15, -6, 10, 5, -1, -1, 0, -7, -6, 4, 17, 12, -6, -2, -11, 3, -6, -4, 0, -15, 3, -15, -9, -17, 13, -16, -13, -15, -15, 0, 0, 1, 10, 4, -5, 12),
    (1, -5, -5, -16, 17, -2, 5, 10, -29, 6, -7, -30, -6, -3, 12, 11, -6, -10, 8, 22, 6, 7, 4, -13, 7, -2, -4, -24, 13, -2, 3, 3, 7, 2, -20, -7, 16, -8, 9, -7, -7, -11, -4, -1, -8, 17, -23, -6, -23, -12, 14, 26, 0, 11, -10, 6, 5, -10, -5, -2, -1, 9, 13, 14, -5, 6, -2, -14, -3, 0, -2, -10, 18, -12, -2, 11, 0, -11, -9, -3, -10, 1, -4, 4, 1, -22, 2, 2, -14, -10, 1, -2, 2, -5, -4, 20, -8, -3, -3, -4, 15, 6, -2, 11, -14, 11, -6, -12, 1, 2, 0, 14, -3, -11, -9, 18, 2, 19, -1, -9, 5, 6, 9, -18, 7, -4, -5, -9, -3, 8, -13, -6, -1, -4, 1, -6, 3, -1, -11, 4, -14, 11, -2, 11, 6, -12, 2, 25, 14, 14, -11, 4, 9, -10, 7, 1, 6, 3, -1, 4, 1, -2, 0, -13, 4, -3, 7, 0, 3, 9, 10, 11, 8, 0, -9, -9, 1, 4, 4, 6, -6, -36, -6, -3, -14, -1, 6, 11, 7, 11, -2, -2, -16, 7, -2, 7, 11, -5, -12, 0, -19, 3, -16, -1, 1, -10, -3, 3, -1, -6, 0, 15, 10, -12, -5, -2, 7, 8, 8, 6, -19, -14, -28, 1, 1, 1, -6, 3, 8, -5, 0, 1, 1, -21, 6, 2, -12, 4, -7, -2, 6, -3, 9, 15, 7, -6, 4, 9, 3, -3, 14, -5, -3, 2, -7, 3, -7, 6, -3, 0, 3, -5, -10, 1, 8, 0, 6, 4, -15, -6, -10, -5, -10, 11, 0, -5, -21, -6, -9, 0, -14, -6, 6, 3, 2, -6, -2, 10, 8),
    (-1, -9, 1, -1, 2, -7, 5, 13, -14, 20, -1, -14, -1, -1, 3, 15, 9, -1, -11, 15, 7, 5, -5, -4, 7, 11, -4, -6, -6, 7, 2, -22, -2, -7, -1, 2, 25, 1, 0, -2, -9, 13, -6, -17, 0, -1, 2, 13, 19, -19, 14, -4, 11, 5, 6, 10, -4, 5, -1, -18, 4, -7, -5, -14, 9, 2, -6, -17, -8, -3, -14, 5, 3, 23, -12, -10, -14, 8, 0, -2, -11, -4, 0, -6, 24, 1, 4, 0, -6, -22, 3, -5, 2, -5, 0, -5, -2, 6, 5, 2, 0, 8, 1, -8, -14, 22, -7, -3, -5, 6, -3, 15, 24, -15, 11, 9, 5, 0, -7, 5, 11, 17, 9, 7, -12, 5, -4, -13, -7, 14, -6, -16, 23, 10, 1, -9, -2, 3, 19, 8, 3, 14, -4, 10, 14, -9, 16, 1, 10, 2, 11, 6, 7, 13, -2, -4, -26, -14, -6, -2, -11, 14, -16, -31, 11, 16, 13, 2, 2, -14, 5, -13, -35, 13, 4, -39, -3, 25, -14, -6, -21, -17, 14, 4, 17, 9, -10, -4, -9, -19, -15, -12, -12, -12, 3, -9, 17, 15, -1, -6, -7, -49, 7, 0, -4, 6, -4, 9, 26, -26, 0, -5, 20, -20, 7, 4, 5, 9, -28, -8, -29, -8, -12, -1, -15, 9, -26, -5, -4, 6, -11, 8, -6, -43, 15, -10, -6, -16, -3, -62, -15, -45, 1, -14, -36, -31, -20, 2, 1, -9, -29, -9, -16, -6, -46, 6, -4, 13, -41, -57, -20, -31, -26, 2, -35, -17, 14, -26, -24, -21, -33, -63, -16, -52, -29, 6, 13, -13, -15, -22, -12, -19, -30, -13, -12, -14, -34, 2, 16),
    (-8, 4, -25, 4, 1, -7, -9, -7, 13, -9, -2, 2, 2, -3, -11, -2, 10, 2, -7, -5, -1, -14, -11, 14, -21, 3, 7, 1, 6, -7, 3, 2, 2, 2, -7, 19, 3, 16, -23, 6, -4, 10, 1, -14, -2, -19, -17, 8, 19, 8, -16, -11, -8, -2, -4, -10, -16, 7, 12, 13, 13, -10, -4, -12, 3, -1, -6, 17, 7, 2, -5, 4, -10, 12, -4, -18, -2, -28, -27, -3, -7, -2, -9, -23, 1, 7, 1, -18, -23, 9, -5, -2, 0, 11, 1, -4, 6, -7, -17, 3, 6, -3, -37, 11, -22, 14, -18, -1, -6, -13, -4, -13, -26, 1, -13, 10, 6, 10, -7, -19, -17, 5, -14, 8, -4, 9, 6, -19, 8, 2, -6, -3, 22, 23, -21, 10, -12, 25, -13, 0, 1, -5, 4, 3, 18, 7, 2, -11, 5, 6, 3, -11, -6, 22, -14, 17, -6, 9, 19, -25, -2, 7, 0, 1, 7, 22, -5, 10, -11, 14, 2, -10, -3, -7, 8, 8, 14, 9, 3, -11, 1, 6, 6, -2, 5, 4, -16, 0, -9, -3, 10, -12, -26, -1, -23, -9, -4, 18, -6, -5, 11, 6, -2, 11, -16, -11, 4, 2, 18, 5, 4, 9, -6, -7, 4, -19, -2, 10, -25, 0, -1, 5, 8, -4, 2, -18, -26, 1, 8, 16, -15, -10, 4, 20, -8, 7, 2, -10, -1, 12, 16, 7, 1, -1, 0, 1, 14, -16, 0, 8, -42, -35, -5, 4, 9, -20, 14, -20, -19, -11, 10, 3, 3, -8, -3, -19, -10, -2, -16, -15, -8, 5, 13, -12, 8, -8, 14, 17, 5, -20, -12, 1, -32, -13, -10, 4, -11, -24, 15),
    (-5, -10, -17, -6, 1, 13, 14, -6, -16, 13, 4, 4, 6, 2, -7, -13, 8, -8, 13, 4, 1, -6, -3, -18, 2, 6, 7, -7, -3, 2, 1, 2, -23, -20, -29, 2, 20, -11, 2, -35, -5, 7, -11, -2, 10, -2, -19, -10, 6, -17, 4, -6, -13, -20, -6, 4, 17, -4, 8, -1, -8, -3, 6, 3, -7, -12, -15, 19, 26, -9, 10, -5, -15, -6, -13, 5, 1, -27, -15, 7, 3, 9, -7, -22, 1, -15, -14, -9, 22, 2, -8, 2, -12, -1, -1, -19, 5, -6, -10, 2, 17, 2, -6, 7, -4, 13, -7, -4, 6, -27, 7, 6, 17, -3, 10, 11, 4, 10, -7, -9, -14, 4, -6, -8, 20, 5, 2, -8, 24, -35, 0, 4, 25, -22, -1, 4, 6, 22, -17, -2, 19, -31, 17, 12, 6, -1, 25, 6, 10, 14, -16, -22, -8, 4, -14, -35, 23, 6, 12, -15, 16, -28, -10, 7, -2, 1, -17, 7, 4, 2, -6, 16, 14, -37, 11, 1, 6, -16, 4, -2, 5, 18, -2, -22, 10, -25, -16, -44, 5, 6, 16, -17, 3, -7, -6, -10, 34, 1, 12, -1, 0, 10, 3, -10, 15, -6, -4, 10, 11, 2, 14, 21, 5, 1, 2, 2, 0, 1, 12, -6, -8, 3, 0, 1, 9, 1, -6, 7, 14, -5, 17, -2, 13, 15, 2, -9, 11, 7, -10, 10, -3, 0, -2, 10, 10, -3, -5, 12, -6, -6, 19, 7, 4, 1, 8, 10, -8, 5, -11, -1, -7, -9, 7, -8, -18, 2, 21, -14, 13, 1, -5, 11, -10, 3, -7, 1, 5, -4, -2, 5, -8, -11, 16, -1, -6, 5, 23, 5, 11),
    (-13, 8, 14, 4, -9, -7, 9, 4, -20, -6, -5, 2, -5, -3, 3, -3, -10, 1, -24, -7, 9, 7, -6, -15, 22, 14, -13, 7, 3, -8, 10, -4, -8, 9, 6, -5, -3, 0, 1, 8, -2, 0, -7, 4, 6, 8, 2, 4, 7, -1, -6, 14, 18, 12, -5, -12, 24, 1, -9, -6, -5, 5, 17, -1, -4, 9, 2, -7, -4, 0, -3, 7, -3, -18, 6, -7, 11, 1, -1, -5, -4, 12, 0, 11, 6, 13, 6, 7, 13, 1, 7, 3, -2, 7, 8, -5, 3, -6, 13, -23, -5, -10, -21, -6, 2, 10, 4, 13, -4, 1, 5, -20, -4, 3, -4, -2, -11, -6, -18, 4, 5, -30, -2, 1, 2, 8, -2, 2, 4, -9, 12, 2, -14, -16, -8, 4, 11, 10, 11, 6, 10, 3, 24, -19, -12, 8, -6, -12, -19, 15, -23, 3, -9, -6, 15, 4, 20, 4, 8, -4, 6, -11, 2, -17, 1, -10, -28, 0, 5, 0, -1, 3, -2, 2, 11, -7, -2, -30, -4, -10, -28, 12, -21, -7, 1, 5, -3, 7, 14, 3, -15, 9, -30, -2, -21, -2, 29, 10, -12, 2, 3, 0, 14, -12, -5, -25, -10, 14, -5, 2, -17, -5, -21, -21, -7, -12, -23, -4, -9, 6, -7, -4, 12, -14, -22, -9, -25, 6, 8, 8, -8, -20, -12, 24, -11, -4, 5, -9, -2, 16, 16, -11, 0, 21, -18, -22, -3, -9, -2, 6, -3, -1, 12, -14, 6, -19, -31, 10, -30, 1, 15, -1, -17, -17, -17, -9, -8, -10, -1, -12, -7, 19, 2, -17, 1, -4, 0, 3, -3, -4, 15, 13, -3, -2, -1, -16, -12, 3, 7),
    (-3, -2, -27, 11, 14, -20, 6, -23, -19, -1, -7, -3, 11, -2, -18, -3, 3, -4, -2, 0, -7, 6, -4, -20, -2, 14, 7, 9, -13, -17, -1, 4, 2, -5, -26, 8, 9, -8, 13, -44, -13, -3, -15, -1, 0, -4, -36, -22, 15, -15, -17, 5, -5, 2, 5, -1, 5, 2, 1, -6, 2, 2, 14, 4, -22, -20, -19, -11, 5, -9, -3, -21, -30, -9, -43, 2, -1, -20, -17, -17, 17, -16, -4, 7, -16, -21, -36, -6, -1, -28, -19, -9, -19, -19, -1, -12, 0, 9, -7, 0, -2, 27, -3, 8, 20, 3, -2, -11, -4, -18, -4, 6, -6, 4, -2, -13, -15, -2, 15, 8, -10, 17, -6, 5, -8, -21, -18, -9, -2, 6, -9, 13, 6, 33, -11, 11, 1, 6, 7, -4, -11, -34, -13, 6, -5, 7, 7, -14, -6, 0, 3, 2, -22, 0, 1, 7, -1, -10, -19, 0, -2, 3, -1, 15, -1, -27, -4, -5, -19, 2, -9, -34, -1, -20, -21, 5, -23, 5, -9, -21, 3, -4, -7, -7, -23, 14, 6, 3, 2, -5, -18, 16, 7, -6, -2, -11, -6, 22, -17, 12, -5, 5, 2, 19, -10, 10, 5, -1, 7, 7, 18, 10, 13, 6, 19, -2, 6, -2, -6, -5, -19, 11, 9, -2, 13, -2, 4, 4, 16, 28, -19, 14, -8, 11, 10, 30, -10, 7, -6, 6, 18, 16, 26, 9, 7, 1, 32, -6, 4, 8, 1, 2, 5, 9, 5, -5, 20, -10, 2, 16, 23, 24, -10, 27, -12, 6, 3, 4, 9, 7, 2, 17, 4, 6, 3, 3, 16, 16, 19, -7, -6, -2, 2, -12, -7, -26, -5, -10, 16),
    (10, 1, 4, -7, -5, -9, 6, -9, 1, -5, 6, -6, 9, -2, -15, 9, -9, 1, 4, 11, -5, -8, 1, 15, 2, 7, 2, -3, -7, 3, 7, 6, 1, 3, -3, -6, 5, 10, 13, 8, 6, -3, 1, -10, -14, -2, -8, -9, -9, 5, 19, 4, 7, -10, 5, 7, -1, 9, 3, 0, 1, 2, -18, 12, -17, -2, -17, 15, 3, 4, -9, 9, 14, 1, -8, -6, -11, -10, 6, -7, 9, -3, -6, -23, -3, 1, -4, -10, 5, -15, -16, 2, 0, -6, -16, 13, 4, -13, 5, 5, -25, -13, 7, 4, 7, 2, 8, -5, 15, 0, 10, -5, -18, 6, -5, 5, -9, 5, -4, 13, -1, -6, 14, -7, 8, 9, -17, 1, 2, -5, 6, 8, 5, 22, 6, 10, -3, 12, -28, 1, -20, -16, 14, 15, -5, -2, 8, 4, -4, 1, 11, -22, 4, 5, 15, -9, 11, 21, -17, -19, 14, -36, -22, 8, 20, 17, -36, 4, -11, -2, -21, 5, -5, -37, -14, -1, 12, -32, 1, -11, 7, 7, 8, -44, 6, -33, -34, -51, -29, -13, -1, -4, -2, -19, 7, 8, -6, -4, 8, 4, -1, 8, -10, 8, 5, 4, 9, 2, -2, -6, 2, -2, -15, 13, 1, 8, -1, 4, 14, 0, 5, 6, 10, -15, -35, -31, 11, -14, -8, 14, -7, -3, -24, 30, -34, 2, -13, -13, 10, -14, 10, -32, 1, 4, -8, 13, 4, -1, 8, -15, 20, 2, -18, 8, 5, -30, -1, -19, -24, -7, 18, 7, 10, -1, 8, -15, -6, -2, 36, -34, -13, -12, -5, -16, 7, 20, -7, 1, -8, -27, -11, -13, -17, -31, -31, 4, -32, -1, 13),
    (-19, -2, -11, -35, 9, -6, 18, -68, 5, 1, 1, 18, 5, -1, -17, -19, -15, -12, -13, -6, -18, -3, -36, -9, -34, -23, 16, 5, -3, -14, 3, 8, -27, -19, -17, -2, 10, -6, 11, -61, -23, 0, 0, 14, 10, -19, -31, -6, -17, -18, -12, 1, 6, -14, -22, -9, -30, 6, 18, -5, -15, -20, 4, 7, -18, -13, 9, 15, -4, -7, 14, -22, -25, 5, -29, 9, -12, -8, -35, 7, 4, -8, -4, 1, 1, -17, -10, -11, -7, 9, -1, -4, -6, -14, -4, -1, 9, 14, -19, -27, 6, 16, 3, -3, -18, 2, 4, -27, -9, -2, -5, 6, -29, 5, 6, 6, 2, 4, -13, 1, -6, -8, 1, 15, -7, -5, 7, -7, 2, 26, -13, -10, 2, 11, 9, 0, 8, -6, 7, -40, -9, 4, -20, -6, -10, 14, -6, -8, -5, -3, -1, -4, -1, -10, 7, 25, 9, 8, 4, 13, -1, 26, 4, 3, -9, -4, 0, 7, 9, -5, 6, -34, -12, -2, -15, 3, 4, 3, -13, -16, -15, -13, 3, -5, -23, 14, 7, 19, 12, -3, -1, 16, -3, 3, -9, 1, 13, 2, -1, 5, -21, -11, -12, 2, 5, -13, -4, 2, 8, -3, 10, 10, -6, -3, 11, -9, -1, 1, -6, -12, -25, 1, -12, -2, 10, 18, 4, 4, -2, 6, 6, 12, 7, -20, -6, 11, 7, 3, 3, -5, 4, 3, 2, -12, -12, -12, 3, -4, 2, 0, -14, 8, 8, 1, -6, 1, 20, -7, 5, 2, 7, 0, -8, 5, 7, -7, -10, 9, 1, 3, 5, -7, 6, -12, 0, -3, -13, 2, -2, -4, -18, 11, -18, -8, 2, -10, -9, -10, 37),
    (-12, 15, 0, -18, -20, -9, 9, -2, 4, -16, 18, 6, 4, 10, -8, -7, -10, -2, -6, 4, -2, -12, -5, 4, 3, -11, 4, 10, -4, -1, -2, 18, -5, -6, 11, -6, -14, -14, -5, -4, 11, -23, 18, 10, -2, 11, -1, -11, -6, -2, -15, 10, 14, -12, 4, 2, 6, -6, -5, 2, 7, -6, 1, 5, -6, -6, 12, 2, -16, -7, -10, 5, -6, -3, 9, -10, 17, 14, 3, -18, -23, -2, -5, 3, 3, -13, -12, -9, 1, -1, -9, -8, 7, -2, 1, 1, -6, -3, -13, 19, 14, 15, -4, 3, 19, 5, -22, -3, -6, -23, 10, 0, -17, 12, -9, -19, 5, 4, 4, -12, -42, -6, -22, -9, 3, 6, 11, 13, 2, 9, -3, 11, -3, -3, 3, 2, 20, 10, -25, -4, -5, -5, 7, 1, -13, 1, -10, -17, -3, 14, 2, -13, -53, -6, 9, 10, 11, 8, 11, 30, 3, 6, 13, 11, -1, -21, 10, -9, 18, 2, -20, 1, 9, -9, -7, 12, -5, 4, -8, -7, -9, 16, 7, -9, -19, 11, 2, 6, 5, 9, 19, 6, -11, 0, 12, 2, -14, -4, -24, -12, -24, -8, 16, -2, 4, 11, -4, 23, 23, -14, -7, 10, 14, -10, 25, -3, 8, 15, -17, -28, -16, -11, -7, -18, -18, -2, 6, -18, 12, 2, -14, -8, -14, -25, 27, 14, 4, 8, -16, 7, 11, -12, 6, -14, 11, -14, 28, 3, 9, 7, -21, -4, -26, -12, -31, 10, -9, -3, 2, -12, 0, 4, -12, 9, 7, -1, 8, 7, -13, 6, -9, -21, -3, -32, 2, -12, 12, -20, -5, 6, 0, -14, -15, 9, -2, -15, -33, 18, -12),
    (4, 15, -9, -7, 14, -2, 2, 0, -5, -4, 2, -1, 4, 3, 9, -11, -6, 10, 2, 3, 1, 3, -11, 11, 0, -8, 12, 5, 1, 3, 7, 2, 0, 17, -10, 7, -12, -12, 15, -4, -17, 7, 14, 3, 10, 21, -1, -14, -2, -2, -13, -6, 10, 1, -2, 9, 3, -4, 6, 14, -15, 0, 22, -2, -14, 13, -13, 10, -6, 4, 8, 1, -13, 4, 5, -4, 5, -6, -3, -18, 3, 0, 0, 3, -2, 3, -2, -9, 13, -15, -6, 12, -7, -12, 4, 5, -5, 9, -9, -4, 1, -9, 9, -6, 0, 2, 2, -16, 21, 2, 1, 8, -15, -3, -5, -9, -18, -11, -4, 10, -11, 12, 9, -14, -6, -10, -41, 15, -12, -7, -10, -15, 1, -21, 0, -6, -3, -6, 3, -10, 17, -2, -5, -4, -8, -6, 1, 2, -12, -11, -20, 10, 1, 5, 7, -22, -7, -6, -28, 14, -12, -1, -5, -25, -2, -21, -3, 7, 4, 9, -4, -19, -14, 6, -8, -15, -18, -3, 1, 4, -21, -21, -34, 0, 11, -8, -5, -6, -2, -2, -6, 8, 17, 10, -14, 2, -6, 12, 3, 11, 3, 8, -3, -11, -15, -10, -9, 9, -6, 5, 4, -9, -14, 9, 7, -15, -12, -8, 5, -5, -3, 8, 6, 2, 15, 6, -13, 13, 8, 19, 13, 20, 2, 2, 7, -14, -6, -17, -9, 14, -17, 23, 18, 2, -23, -8, 6, -8, -16, -22, -21, -2, 2, 6, 8, 2, -5, -7, -15, 0, 11, 10, 10, 15, -18, 28, -10, -20, -9, -12, 1, 19, 0, -18, -3, 6, -18, -10, 10, 7, 1, -21, -5, 2, -8, -20, 9, 5, 4),
    (-7, 9, -2, -2, -5, -9, -10, 11, 12, -10, 11, -2, 11, -10, -10, -4, 12, 5, -1, 6, -10, -1, -13, 5, 4, 12, 6, 15, -10, -1, -17, -13, -18, 19, -2, 7, -2, 0, -1, 19, 1, -10, -1, -14, 23, -12, 12, -15, 6, 18, -29, 8, -6, -6, -7, 6, 10, 14, -6, -1, -14, 8, -18, -27, -3, 15, 6, 1, -6, 6, 2, 19, -2, 1, -5, -27, 8, -8, 13, -13, -18, 11, -13, 3, 0, -5, -2, 2, 17, 6, -11, 1, -16, 1, -12, -7, -3, 1, -3, 7, 19, 10, -1, 7, 2, 25, -11, 6, 9, -1, 20, 11, 21, 2, -11, 5, -11, 11, -14, 7, 6, 2, 6, -8, -7, 3, -7, -30, 10, -1, -7, 13, -6, -4, -7, -1, -10, 15, -3, -1, -6, -1, 26, 15, 13, -26, -14, -1, -10, 26, -4, 9, 4, -4, 3, -10, -7, 7, 19, -27, 11, -6, -9, -11, -2, -4, -31, -14, -5, 1, 0, 4, 7, 6, 5, 4, 3, -32, 4, -11, 15, -8, -5, -3, 5, -16, 12, -3, -6, 13, 20, 1, -12, -3, -26, -10, -5, 9, -21, 0, 0, -11, 10, 4, -37, -1, -2, 1, 19, -5, 1, -7, -23, -15, 14, 4, 4, 8, 0, 11, -9, -3, -1, 9, 2, 6, -22, -17, 10, 1, -3, -17, 1, -25, 11, -3, -16, -17, -29, -24, -2, -10, 16, -2, -14, -31, 15, 1, 3, 11, -31, 19, -3, 2, -30, 2, 4, -16, 1, -33, 3, -9, -13, -6, 14, -33, 0, 4, -2, -17, -16, -30, -8, -14, 17, -4, 14, -10, 12, -28, -8, -2, -42, -16, -13, -6, -8, -3, 23),
    (13, -1, -19, -10, -5, 2, 12, 10, 6, 2, 0, 3, 5, -4, 7, -9, -15, 6, 5, -3, -3, 2, -5, -1, -9, -18, 22, 2, -7, 10, 7, -2, 19, 25, -15, -26, 2, 1, 2, -2, 13, 0, -5, -6, -18, -2, -2, -3, -23, -1, 3, 4, -4, 19, -22, 2, -18, -32, 0, 23, -7, 27, 3, 1, 2, 19, -3, -15, 13, 0, 13, -1, 19, -21, -3, 2, -7, -1, -22, -6, 1, 1, 6, 7, -7, 2, -4, -8, -18, -4, 10, 15, -10, 23, 11, -6, -2, 18, -35, -2, -2, -4, -17, 6, 9, 3, 12, -10, -1, -16, -7, 0, -6, 4, 10, 3, -6, -2, -14, -19, -3, 9, 5, 7, 2, -4, 1, 0, 11, 6, -21, -9, -5, 14, -24, 13, -4, 9, -10, 6, -16, -6, -4, 12, -3, 9, 3, 27, 9, 6, -15, -4, -3, -10, -19, 8, -1, 8, -1, 6, 6, 2, -17, -22, 9, 6, 13, 2, -4, -5, 1, 5, -1, 1, -6, 11, 20, 17, 3, 1, -11, 13, -4, -10, 4, -11, -4, 10, 0, -1, -10, -9, -18, 0, -27, 0, -36, -5, -23, -7, -4, -12, -15, -10, -13, -17, -18, -2, -23, -9, 6, -23, -24, -3, -11, -12, -20, -16, 5, 13, -17, -12, 9, -6, -16, 6, -9, 16, -31, 4, -17, 6, 3, 8, -9, -6, -20, -6, -4, 4, 6, -1, 9, 6, -8, -14, -1, -8, -3, 3, 4, -4, -15, -7, -7, 7, 8, -20, -6, 4, 4, 14, 10, 6, 10, -2, 5, 3, -8, -1, 4, 12, 14, -17, 13, 4, 6, 10, 1, -4, 7, 8, -12, -13, -6, 4, 5, -2, 19),
    (19, -5, -7, -13, 0, 14, 3, -3, 6, -5, 10, 2, -14, -4, -22, 1, -4, -5, 20, -7, 1, -5, 0, -5, -6, 2, -1, 4, 4, -15, 7, -6, 6, -2, 12, 18, -13, 3, -6, -2, -7, -4, 16, 0, -8, -6, -3, -8, -11, 9, -10, -14, -8, -7, 4, 5, -3, -14, 1, -2, 16, -11, -10, 30, 19, 3, 6, 1, -8, 8, -6, 9, 22, -2, -8, -5, 9, -6, -21, 8, -6, 2, -7, -10, 5, -3, 2, -5, -6, 15, -4, -4, 19, -6, 3, 11, -9, 7, -1, -25, -8, -13, -6, 12, 15, -7, 6, -7, 3, 10, -8, -8, -11, 11, -3, -1, -24, -6, -24, 4, -2, -10, -14, -6, -16, 1, 8, 6, -2, -7, 10, -11, -10, -1, -26, 9, 12, -19, 17, 13, -9, 17, 6, -10, -6, 14, 10, -5, -17, -7, -9, -2, 1, -7, -41, 21, 6, 10, 14, 21, 11, -9, 14, -9, -9, 13, -2, 12, 10, 4, -3, 17, 17, 17, 19, 13, -6, -14, -2, 3, 1, -24, -9, -3, 4, 1, -25, -1, 11, 6, 7, 9, -19, -2, -43, -13, -8, 0, -7, 1, 6, 14, 3, -19, 12, -22, -6, 15, -11, -6, -12, 7, 0, 9, -7, -28, -20, 0, -9, -17, -3, 3, -7, -44, 1, -5, -8, -3, 0, -12, 0, -1, 10, 11, -44, -21, 11, -29, 3, 18, -13, 3, 0, 14, 17, 26, -14, -17, -10, -21, -4, -18, 14, 4, 3, -37, -25, -17, -7, 6, -19, -12, -20, -15, 15, 2, -20, -17, -16, -16, -4, 6, -25, -10, -5, -6, 2, 1, -14, -22, -18, -24, 7, -11, -1, 4, 12, -37, 2),
    (19, -16, 9, 22, 16, 5, -4, 15, -3, 19, -7, -16, 7, -20, 4, 28, -7, 0, 12, 6, 15, 12, -3, -2, -5, 13, -24, -18, 10, 11, -1, -23, 26, -42, -15, 16, 14, -2, -25, 12, 1, 22, -19, -31, -5, -51, 9, 22, -1, 8, 19, 5, 12, 21, -7, -24, -6, 1, -23, -42, 28, 6, 5, -39, 4, -19, -27, 0, -8, 2, -15, 4, 7, -10, -12, -3, 5, -38, 5, -12, 4, -8, -6, -21, -16, 13, -5, -31, -1, -22, -7, -16, -1, 2, -6, -34, 10, -13, 10, 9, 5, 2, -7, -2, 18, 10, -2, -7, 11, -9, -6, 14, -11, -2, 22, 9, 2, 4, 6, 8, 0, 18, -6, -9, 0, 4, 2, 2, 7, -20, -3, 15, 6, 5, -10, -2, 8, 7, -1, 5, 1, -10, -5, 14, -10, -13, 16, 11, 15, 4, 7, 11, 4, 7, 6, -8, -7, 4, 2, 6, -5, -10, -13, 2, -14, -1, 0, -3, -21, -7, 2, 2, 14, 4, 3, -30, 4, -9, 9, -3, 6, -6, 3, -12, -1, -4, 6, -3, -12, -3, 0, -3, 9, -14, 10, 1, -1, -1, 7, -8, 6, -4, 8, -1, -3, -1, -7, 0, -5, 0, 2, 1, -11, -9, 3, 1, -3, 2, 0, 1, -1, -12, -7, 2, -1, -13, 8, -1, 3, 4, 10, -4, -1, 0, -2, 8, -2, -3, -13, 2, 5, 11, 8, 6, 7, -22, 17, 0, 2, -2, -6, -11, -7, -2, -2, -6, 6, 5, -4, 14, -3, 8, 7, 5, -4, -14, 5, -8, 5, -3, -10, 11, -6, 9, 6, -10, 12, 4, 5, -13, 0, -22, -16, -8, -9, -4, 9, -7, 16),
    (2, -17, -18, 5, 1, 20, -5, -4, -6, 14, -8, -10, 23, 2, 1, -5, -17, -7, 6, 5, 2, -2, 8, -13, 0, 11, -4, -16, 0, -7, 7, -21, -17, -57, -19, 14, -3, 16, 1, -3, -11, 0, 2, -1, -9, -2, -23, -3, -3, -19, 3, -21, 4, 12, 19, -7, -4, 2, -2, -14, -2, -26, 8, 8, -13, -23, -9, -10, -14, 9, 4, -6, 8, -2, -21, -10, -12, -36, -23, 9, -16, -20, 12, -21, -10, 12, -4, -7, -5, -26, -2, -4, 7, -32, -3, -17, 17, 3, -17, -8, -9, 0, 11, -2, -1, 0, 3, -12, -8, -4, 12, 5, 4, -5, 9, -3, -4, -2, -19, 1, -35, -12, 5, 11, -7, 8, -9, 14, 11, 3, -15, -19, -2, -2, 2, -6, 4, -21, 7, -34, -5, -11, -17, -7, 2, 7, 13, 9, 6, -6, -1, 0, -30, -8, 0, 22, -4, 20, -15, 38, 1, 12, 2, -14, -23, -6, 6, 7, -13, -10, 4, -21, 3, -2, -17, -18, -15, 3, 5, 7, -10, -24, -1, 7, -6, 0, 11, 2, -5, 8, -15, 15, 16, -17, -29, -13, 4, -2, -19, 7, 14, 4, -7, 3, 0, -11, -13, -8, -14, 11, 6, 8, -5, 15, -7, -9, -6, -22, -16, -4, -6, 17, 15, -21, 5, -5, 5, 1, -8, 5, 5, 22, 19, 4, -10, 6, 2, 1, 20, -5, -18, 18, 7, -2, -15, 15, -2, -13, -2, -12, -13, -3, 14, 21, 14, -18, 5, -22, 11, 9, -1, 0, 15, 13, -6, 6, -12, 11, -8, -2, 18, 6, -1, -9, -8, 6, 0, 5, 2, -3, 6, 14, 12, -7, 9, 11, 14, -13, 9),
    (2, 0, -10, -18, -2, 2, 10, -2, -21, -1, -10, -13, 9, 7, 7, -1, -5, -27, 8, 30, 8, 19, -14, -6, 8, -15, -25, -10, -1, 4, 19, -19, 3, 10, -19, -23, 9, -23, 11, -20, -4, -25, 6, -5, -13, 2, 13, -2, 2, 0, -4, 18, -4, -14, -10, 12, 3, -26, 16, 1, 8, 15, 4, -9, 6, -7, -29, -13, 1, -17, -19, -14, 2, -9, 10, 7, -24, -29, -33, -16, 3, -21, -6, -10, -9, -4, -8, -17, -5, -2, -2, -10, 4, -23, 2, -8, -7, 0, -4, -16, 5, -6, 3, -6, -5, 2, -1, 6, 2, 10, 3, 4, -11, -12, 0, 15, 7, 14, -11, 0, 13, -11, 4, -9, 1, 11, 14, 8, -5, 12, -10, -10, 18, -2, 26, -10, 13, 4, 7, 7, 10, 0, -9, -21, -26, -1, 2, 10, 13, 14, -6, -10, 13, -5, 4, 5, 2, 6, 25, 4, -9, 11, -1, -3, 3, 6, 14, -5, 7, -8, -7, 3, 3, 4, -9, -3, 0, 5, 6, 11, 11, 17, -2, 3, 15, -6, 7, -2, -13, 8, 17, -22, 8, 6, -8, 1, 15, -2, 7, -4, 4, 2, 11, 0, 5, 1, 2, -2, -7, 8, 3, -5, 16, 6, 3, 2, 1, 1, -13, -4, 0, 2, 1, 1, -2, 10, -1, 6, 0, -11, 11, -8, 12, 12, -1, -9, 19, -3, 2, -1, -2, 1, -2, -2, 20, 12, -18, -2, 6, 2, 9, 16, 6, 1, 10, -3, -18, 2, -2, 1, 5, -9, -5, 0, 0, -2, 8, -10, -1, -5, 6, -17, -3, 1, -14, 10, -9, 12, -14, 2, 4, -12, 5, 1, 6, 8, -9, -3, 5),
    (-11, 4, -1, 10, -12, 4, -7, -13, -10, -8, 7, 1, -8, -10, 0, 8, 15, -6, 13, -7, -8, -20, 9, -14, 11, 21, 1, 10, -15, -15, -17, 6, -13, 2, -3, 29, -14, 11, -7, -3, 3, -15, 2, 0, 3, 2, -1, 10, 22, -6, 1, -3, 1, -13, 15, -15, 19, 22, -12, 13, -20, -2, -11, 11, -10, -8, -4, 7, 8, 6, 2, -16, 4, -10, -11, -2, 10, -3, 2, -4, 1, 4, 2, 5, 3, -6, 8, -6, 2, 17, -10, -5, -2, -7, -18, 2, -8, -7, 12, 4, -2, 10, 11, -22, -18, -7, 22, 2, 8, -7, -27, 5, 12, -3, 2, -42, -5, -30, 6, 13, -6, 14, 16, 11, -4, -26, -3, -5, -19, 2, 18, 14, -4, -7, 4, -14, -20, -1, 10, -3, 13, 6, -17, 1, 9, -16, -8, -7, 3, 0, 14, 10, 5, 19, 19, -3, -17, -15, -21, 4, -9, 5, 10, 14, 5, -5, -1, 3, -3, -8, 5, -7, 2, 5, 2, 13, 13, -7, -11, -1, 5, 5, 4, -10, 10, 4, 8, -7, -6, 1, -39, 11, 14, -17, -11, -15, -4, -3, 12, -34, -2, -12, -12, 1, -8, -11, -13, -3, 10, -6, 8, 8, -9, -15, 3, 2, -3, 4, 9, -4, 0, -19, 0, -1, -11, -9, -5, -22, 13, 10, 7, -6, 2, -10, 10, -15, -17, -15, -7, -11, 3, -9, 14, 12, -6, -15, 3, 4, 3, 7, -5, 13, -5, -15, -10, 4, -12, -6, 8, -9, 5, 2, 4, 9, 14, -1, 0, 0, 0, -6, -2, 2, -5, 2, 15, 1, -5, 15, 1, -2, 9, -8, -8, 5, 6, -9, 7, 5, -4),
    (5, 7, 2, -3, 14, -19, 16, 2, -11, 9, 8, -10, -15, 11, 13, 17, -4, -13, -8, 11, 6, 9, -26, 18, -2, 5, 10, 9, 5, 0, 2, -10, 10, -6, -10, -4, 8, -15, 11, -6, -14, 14, 4, -5, -3, 6, -6, 25, -3, -5, 2, 20, 19, 14, -3, -11, -5, -1, 17, -3, -6, 8, 7, 0, -7, -3, 3, -3, 12, 3, -3, -10, -15, -2, -10, 1, -7, 5, -14, 3, -5, -13, 17, 7, 7, 7, -1, -3, -9, -13, 7, -2, 3, -1, 1, 4, -17, 6, -14, 11, 2, 4, -21, 0, -2, 6, -9, -15, -12, -15, -11, -6, 6, -16, -2, -14, -17, 2, 2, 9, 3, 26, -2, 1, -6, 5, -41, -16, -11, 13, -8, -2, 18, 1, -9, 10, -4, 6, -6, -17, -16, -8, -6, 19, -3, -16, 10, 12, 5, 2, 3, -6, 0, 18, 8, -14, 5, 14, -5, -7, -3, 5, -10, -10, 6, -8, 0, 0, -2, -8, 2, -16, -2, -4, 0, 15, 6, 4, 5, 6, 2, 13, -9, -2, 0, -15, -5, 7, -2, -1, -8, 3, -3, 10, -7, 6, 11, -23, -6, -15, -5, -11, -26, 1, 5, -28, -9, -19, -11, 4, 2, 0, -39, -5, 12, -3, -7, 8, -1, -13, -11, -22, -36, 5, -22, -25, 15, 15, -6, 0, 4, -8, 2, 12, 7, 2, 17, -2, -16, 3, -3, -2, 10, 3, -4, -19, 2, 7, 1, 11, -18, -27, 10, -10, -16, 5, 10, -11, -9, -13, 15, 10, 2, 15, 2, 11, -2, -2, -1, -3, 3, 10, 6, -22, 20, 13, 2, -4, 8, -3, 9, 4, 10, -19, 0, -6, -4, -6, 16),
    (-14, -8, 17, 24, -1, 0, -18, 17, -16, 1, -18, -9, 3, 2, 1, 6, 14, -10, 1, 8, 7, -6, 13, -11, 11, 8, -16, -12, 6, -11, -6, 6, -8, -19, 8, 10, -2, -6, -8, 7, -30, -3, -11, -4, 2, 8, 4, -5, 9, 6, -2, 3, 11, 10, 12, -9, 8, 9, -1, -3, -16, -9, 4, -3, 16, -10, -9, 2, 2, 10, -6, -1, -11, 1, 3, 3, 5, -6, -12, 9, 5, 5, -6, 7, -10, 1, -8, -6, 4, 1, -1, 0, -23, 3, -2, -10, -19, -9, 12, 22, -15, 6, -8, 10, -17, 6, -11, 12, -2, 3, 26, -6, 1, -20, -20, 10, 2, 9, 10, -9, 17, 11, -1, -18, -1, -1, -17, -5, -9, -7, 6, 15, -8, 21, -2, 9, -8, -5, -17, 14, -16, 2, 14, 0, 6, 1, -10, 22, 8, 20, 10, -3, 19, 15, -1, -16, -14, -5, 3, -6, 8, -7, -7, 14, 5, -1, -9, 6, -21, -4, -1, -14, 9, -1, 3, 16, 7, 4, -5, 16, -9, 13, 2, 1, 10, 1, -7, -2, -14, -6, -6, -9, -5, -9, -2, 1, 6, 4, 4, 6, -7, 16, -17, 8, 6, 2, 11, -7, 1, 13, -4, 4, 1, 18, 4, 0, 1, -13, 1, 3, -3, -3, -3, -12, -5, 5, 3, 10, -5, 3, -2, 1, -7, -1, -4, 8, -2, 5, 13, -1, 0, 10, -5, 8, 6, 23, -5, -4, 5, -11, 9, -2, -14, 2, 15, -1, 13, -2, -3, -28, 1, -9, 5, -11, -7, -2, 2, 2, -1, 4, 5, 7, -1, 6, -2, 12, 23, -6, 4, 1, 6, -21, 12, -6, -11, -5, 1, -11, -10),
    (11, -17, -29, -19, 0, -14, 18, -25, 5, -2, -2, -4, -22, -4, -6, -14, 2, -17, 8, 6, 5, 10, 0, -8, -16, -18, 7, 2, 11, -8, 13, 15, 7, 4, -12, -12, -15, -12, -7, -22, -2, -15, 9, 13, 0, 8, -44, 0, -1, -6, 11, 2, 16, 6, 1, -12, -20, -17, 5, 22, -1, 2, 11, 3, -5, 4, -13, -4, -3, 7, 8, 3, 10, -10, 10, 5, 9, 8, -43, -4, -5, 11, 2, 6, 10, 8, -6, 7, -4, 5, 6, 13, -21, 6, 0, 2, 5, 9, 2, 1, -6, -7, -20, 2, 12, -12, 2, -7, 5, -17, -21, -24, -22, 9, 12, -17, -9, -4, -5, -2, -3, -1, 6, -2, -3, 1, -27, 23, 1, -3, 17, 9, -19, -5, 2, 16, 21, -6, 6, 8, 18, 2, 6, -21, -28, 2, -20, 4, -17, 5, -9, -5, 1, 0, 14, -10, 11, 5, -26, -2, -3, -3, 10, -2, -13, 8, -10, 10, 2, -9, -11, -13, -7, 1, 15, -10, -6, -8, -16, 0, -20, 16, -1, -10, 6, 5, -6, -17, 8, -1, -12, -11, -25, -23, -13, -16, 17, 14, -5, 7, -2, 7, -7, -1, 4, -7, 10, 10, 8, 6, -10, 2, 5, -10, -5, -1, -8, -9, -2, -5, 3, 2, 7, -17, -26, 1, -31, 1, 4, 18, -4, -1, 0, 18, -6, 7, 6, -10, -2, 11, 3, 2, -10, 3, 12, -3, -3, 7, -2, -4, 1, -1, 10, -12, 13, -5, -13, -7, -19, -11, 10, -7, -5, -15, -3, 21, 10, -14, 10, -3, -10, 19, 11, -4, -2, -3, -13, -12, -2, 12, 2, 1, 7, 12, 3, -20, 11, 10, 33),
    (7, 18, -5, -6, 5, -10, 8, 3, -24, -6, 2, 12, -1, -14, -4, -2, -16, -2, 0, -1, -5, 0, -4, -2, -20, 0, 10, -2, -5, 15, 2, -4, 20, 3, -13, 0, 15, -12, 23, 3, -9, -5, 8, 2, -2, -2, -15, -2, 3, -7, -6, 0, -9, -2, -10, -9, -38, -6, 2, 19, -21, 21, 15, -8, 13, -5, -14, -5, 1, -1, 7, -1, -5, -3, 5, 8, 12, -10, -22, 4, -26, -3, 6, -5, 3, -4, -4, -9, -14, 21, -1, -2, -10, 10, 20, -3, -19, 0, 10, -6, 5, 14, -4, 5, -16, 3, -25, 1, 4, -23, 6, 10, 10, -12, -3, 2, -11, 4, 6, -9, 3, 3, 13, -1, 9, 0, -11, -26, 10, 10, -16, 8, 14, 14, -38, 11, 22, 6, -18, -14, -14, -23, 1, 5, 13, 1, 18, 5, -2, 8, -9, -10, -10, 4, -29, -4, -1, 10, 7, -13, 25, 13, -22, -1, 4, -6, 9, 14, 20, -5, 1, -21, -17, -10, -9, 30, 9, 22, 6, 5, 0, -1, -21, -7, -22, 40, -16, 7, 12, 17, 13, 15, -16, -16, 6, -20, 5, 2, -5, -33, -34, 7, -7, 3, 7, -15, 2, 2, 13, 12, -8, 12, -9, -21, 2, -6, -7, 5, 17, 9, 14, -16, 6, -29, -19, -12, -28, -14, 4, 11, -10, -4, 4, 8, -21, 10, 18, -22, -14, -8, 4, 1, 1, 7, -5, -24, 2, -6, -1, -6, -24, -25, -6, -5, 7, -18, -3, -24, -27, 17, 2, 5, -10, 2, 7, -7, -25, 1, -16, -22, -5, 10, 0, -11, 12, 7, -6, -4, -17, -15, -10, 20, -30, -9, 5, 8, -6, -22, 4),
    (-30, -20, 0, -13, -1, -6, -3, -19, 0, -14, -20, 5, -6, -30, -1, 5, 1, 7, -13, -16, -23, 3, 3, -5, -25, 20, -2, -32, -2, -11, -6, 7, -55, -14, 6, 11, -15, -17, -3, -5, 22, -19, -35, 2, 2, -26, -2, -12, -2, 12, -11, -30, -7, -6, 3, 6, -23, 9, -33, -3, 13, 18, -3, 27, -50, -12, -14, 35, -5, -3, -12, -5, 11, -3, -26, 1, -31, -15, 10, -4, 1, 1, -19, -23, -7, -31, -7, 10, 11, 15, -18, 2, 6, 6, -2, 12, 14, -17, -7, -9, 1, -2, 5, 0, -26, 8, -1, 13, -20, 10, -5, 19, -43, 1, 8, -2, 10, 6, -14, -2, -3, -6, 3, 3, -6, 5, 14, -11, 23, -11, 2, -4, 4, -22, 2, -14, -40, 3, -1, -19, -26, 20, 11, 11, -27, -6, 7, -3, 14, 6, -6, -8, -12, -27, 1, 14, -15, 4, 34, -1, 9, -10, 15, 10, 13, -32, 0, -18, -26, 13, 0, 17, 5, 18, -3, 7, -8, -14, -17, -6, 23, 3, 0, -6, -21, -8, 19, 5, -6, 2, 31, -8, -14, 12, -13, 1, 9, 8, -11, 15, 14, 2, 6, -7, -8, -14, -2, 12, -4, -18, 10, -2, -2, -3, -5, -2, -5, 13, -12, -1, 7, 10, -17, 4, -15, 17, -22, 0, 13, 9, -12, 9, 18, -9, 10, -11, -14, -19, -13, 14, 6, -11, 16, 7, 6, -11, -8, 1, -5, 11, 5, 16, 2, 10, -15, 8, -15, 14, -17, 21, 10, 10, -25, 6, 21, -1, -1, -12, -34, -12, -8, 3, -6, 20, 5, -9, 0, -8, -9, 6, 0, -6, -16, 14, 8, -2, -6, 16, 1),
    (1, -8, -10, 14, 24, 2, 6, -7, -11, 15, 2, -5, -9, 2, 2, 14, 7, -15, 15, 1, 8, 10, 8, -2, -4, 5, 9, -2, -4, -2, 8, -2, -1, 13, -8, 11, 22, 2, 6, -2, 9, 8, -7, 11, -18, 6, -25, -6, -8, -11, -3, -19, 14, 15, 4, -28, -33, 2, 5, 13, -1, 9, 10, 10, 0, 2, 9, 12, -38, -18, 3, -2, -22, 5, -6, -3, 5, -2, -16, 8, -11, -1, -12, -10, 9, 4, -2, -23, -15, 10, 2, 3, -5, 2, 7, -3, -5, 15, -2, 8, 9, 10, -18, -2, 15, -11, 2, -5, -16, 2, -10, 17, 11, -13, 22, -10, 18, -6, 12, -12, 0, 4, 2, 12, 4, 4, -11, 15, 1, 21, 2, 5, 7, 7, -8, -3, 19, -10, 17, 5, -12, -2, -22, 10, 8, 7, 12, -10, 19, -1, 8, -17, 7, 0, -16, 17, 9, 2, -25, 18, 4, 8, 6, 1, 5, 7, -7, 4, 13, -5, -1, -2, 6, -3, -10, 2, 16, 6, 12, -10, 4, 5, 2, -16, 5, 37, -10, -4, 10, -5, -12, 10, 2, -11, 21, 2, -16, -6, 5, 4, -1, -13, -14, 2, 1, -7, -10, -9, -12, -7, -4, -19, -20, -3, 1, -8, -6, 11, -2, -15, -2, -7, -20, 15, 11, -27, -9, 13, 0, -11, 21, -16, 2, -9, -23, 0, 2, -22, 1, -21, -13, -3, -2, -14, -32, 2, -6, -1, -10, 10, -19, -36, -2, -13, -7, 16, 11, -21, -27, 11, -1, -28, -13, -28, 12, -5, -56, -3, -3, -13, 5, -16, 6, -16, 3, -6, 0, 8, -12, -2, -5, 37, -11, -16, 0, -14, -2, 5, 17),
    (5, -9, -1, 11, -4, 15, 5, 1, -27, 8, -2, 3, 0, -4, -10, 11, 8, 14, 4, 1, 1, -4, 0, 5, -6, -1, 4, 7, 16, -2, 14, -7, -5, -4, -5, -4, 5, 0, 1, -1, -15, 7, 8, -2, 8, 10, 10, 15, 10, 2, 1, 10, 7, 2, -2, 13, -4, -16, -2, -18, -3, -10, 7, -7, -7, -1, 2, -6, 4, -5, 2, 2, -14, 0, 11, -4, -8, 3, -2, -1, -8, -12, 3, 1, -1, 9, -2, 3, -6, -20, -15, -13, 0, -5, -4, 0, 3, -10, -12, -27, -8, -5, 8, -12, -9, -10, 7, -11, 3, 7, -38, -10, 3, 10, 0, -39, -5, -22, -4, 20, -6, -7, -8, -11, -2, -3, -1, 10, 0, 7, -8, -21, 1, -17, 3, -8, -13, 4, 16, -26, -5, 7, -8, 0, -6, 5, 6, -4, 6, -19, -3, 24, -8, -22, 6, 0, -5, -7, -11, 4, -2, 2, -6, -8, 10, -11, -2, -8, -23, 12, 6, -9, 9, 6, 3, -8, -18, -6, 7, 2, 2, 8, -1, 12, -14, -20, 2, -1, -9, -6, -23, 15, -5, -6, -4, -1, 9, 5, -3, -2, 5, -15, 5, 3, -1, -6, -1, -3, 6, 3, 2, 1, 6, -19, 0, -1, 0, 2, -11, -6, -6, 0, -7, 10, 2, -4, -15, -1, 18, -8, 11, -2, 0, -15, 4, -8, 12, 10, -6, -5, -3, -5, -5, 0, 0, -14, -4, 5, 2, 7, -7, 10, 17, -6, 1, -2, -11, 8, 1, 3, 7, 16, -3, 2, 8, 12, 10, -9, -1, -1, 0, 8, -2, -6, 2, 5, 4, -6, 14, 8, -4, -2, 8, 11, 9, -2, -8, 4, 19),
    (-3, 4, 4, 10, 11, 8, 2, -2, -8, 8, -26, -8, -17, -10, 17, 7, 6, -12, -21, 16, 5, 3, 4, -7, 4, 2, -1, -5, 4, 1, -4, -28, 10, -28, -47, -5, 10, -22, -19, -14, -9, 5, -27, -4, 2, -26, -11, -8, -7, -17, -15, 18, -13, 9, -23, -5, -8, 0, -25, -13, -10, 12, -10, -37, 3, -28, -36, -8, -5, -6, 1, -7, -8, -6, -19, 2, 5, -18, -3, -18, -15, -9, -13, 10, -22, 4, -13, -11, 11, -7, -20, -7, 1, 3, 2, -12, -1, 8, -1, 3, 8, 29, -9, 11, -16, 6, -2, 11, -13, -14, 5, 3, 41, 2, -10, 9, 7, 6, 9, -34, 18, 19, -3, 6, -1, 5, -2, -8, -6, -2, -11, 0, 24, 14, 2, 1, -11, -4, 0, -29, -16, -7, 2, -2, 17, -5, -6, 3, 9, 7, 10, -34, 7, 6, 14, -4, -21, 5, 10, -10, -4, 6, -3, -6, 5, 4, -6, -10, -24, 0, 0, 5, 9, -3, -6, 8, 17, -8, 12, 5, 0, 0, 9, -25, -3, 20, 6, -5, -8, 3, 13, -7, -30, -12, 4, 10, 13, 4, -22, -5, -5, 1, 4, 7, -10, -1, 2, 7, 10, -2, -14, -5, 30, 6, 5, -13, 12, 6, 8, -1, -5, 2, -7, 11, -24, -3, 7, 25, -6, -3, -18, -5, 17, -3, 0, 11, -2, 0, -2, -2, 14, 9, -11, -20, 25, 5, 1, -5, 10, 14, -3, 14, 10, 6, 7, 12, 6, -16, 5, -7, 6, -7, -9, 3, 14, -10, 8, 8, 8, 2, 5, 13, 8, -13, -7, 1, 22, 10, -5, -2, 2, 15, 2, 11, 8, 5, 21, 4, -9),
    (-18, 14, -8, -11, 10, 3, -2, 6, 1, 3, -2, 3, 4, -4, 3, -9, -1, -2, -2, -2, 0, -1, 6, 10, -6, -15, 0, 1, -8, -18, -17, -1, -22, 20, -19, 2, 16, 10, -3, 9, -14, 3, 6, -3, 9, -12, -1, 8, 22, 2, -5, -6, -5, 3, 5, 10, -5, 7, 1, 12, -15, -14, -14, 1, -12, 9, -10, -9, 12, 10, 3, 4, -3, 3, 4, -6, -4, -19, -8, 6, 10, 10, -2, 0, -17, -3, -6, 8, -3, 16, -6, 14, -10, -13, -21, 1, 9, 7, 6, -22, -21, 8, -13, -4, 11, -2, 6, 22, -13, 15, -7, 3, 12, -17, 3, -7, -3, -8, 16, -6, 22, -4, -17, 4, -4, -10, -13, 16, 15, -3, 10, -4, -2, 11, -18, 5, 0, -6, 14, 32, -9, 8, 2, -2, 12, -11, 1, 2, 6, -4, 28, -2, 15, -14, -11, 1, 15, -2, -9, 6, 14, -6, 1, -5, -4, 5, -26, 12, -8, -4, 10, -2, -14, -10, 4, -10, 4, -12, -10, 1, -3, -8, -2, -16, -19, -24, 3, 2, 11, 4, -5, -6, -2, 1, -20, 5, -20, -7, 9, -3, 3, 3, -25, -7, 10, -30, -1, -8, -11, -3, 0, -8, -22, 4, -12, -6, -31, -9, 5, -18, -9, 1, 0, -8, 4, -7, -7, 13, -22, -7, -15, -5, 11, 19, -17, -6, 0, -42, 0, -3, -14, 8, 2, -11, -15, 10, -5, -16, -26, -19, -3, 1, 14, 4, 21, -6, -9, -21, 0, 7, -5, -12, -15, -8, 1, 0, -12, -1, 19, -19, -11, -11, 2, 24, -2, 8, -2, -17, 2, -17, 5, 12, 2, -8, -1, 10, 22, -19, 18),
    (34, 18, -18, -11, -9, 18, 10, 11, 17, -1, 16, -9, -21, -13, -18, -14, -18, 15, -2, -25, -12, -3, -15, 4, -34, -19, 12, 16, -7, 14, -8, 9, 16, 16, -9, 6, -18, 13, -5, 15, 9, 1, 15, -17, -12, 5, -16, -6, -8, 9, -15, -19, -19, -24, 3, 4, -30, -18, 13, 14, -17, -7, -18, -2, -1, 12, 6, 8, -15, -22, -6, 10, -6, 14, 12, -17, -7, 2, 2, 8, 15, 7, -10, -4, -9, -17, 13, 5, -12, -9, 2, 6, -1, -10, -22, 5, 5, -1, -8, -15, 0, 22, -31, 17, 13, -10, -13, 18, -12, 2, 8, -3, 33, 0, 7, -2, -14, -9, 11, -7, -6, -2, -26, -22, -18, 22, -6, -10, 0, 11, -14, 0, 8, 23, -9, 26, -7, -18, -3, 25, 6, 6, 7, -5, 22, 15, 4, -6, -14, -9, 5, 2, -5, -5, -10, -2, -10, 2, 4, -10, -6, 5, 5, 8, -1, 13, -14, 7, -3, 17, -2, 12, -6, 2, 4, -3, -3, 6, 8, -2, -11, -6, 10, 3, -11, -7, -10, -3, -5, -12, -14, -2, -4, -8, -4, -7, -2, 1, -8, -18, -3, -1, -9, 10, -8, -9, -1, 1, 5, -4, -15, -1, -6, -7, -2, -4, -3, 2, -4, -11, -20, -8, -14, -3, -5, -25, -5, 2, -1, 6, -15, -7, 3, -11, 1, 17, -7, 7, 0, 6, 14, -1, -4, 8, 25, 1, -12, -4, -1, 6, 3, 5, -2, 10, 2, 0, 0, -11, -6, -13, -6, 0, -14, -16, -1, -10, 11, 12, 6, 12, 4, 10, 6, 14, 1, -1, 2, -1, -2, 6, -2, -2, 14, 4, 1, -2, 11, 5, 17),
    (17, -28, 13, 2, 11, -3, 18, 6, -8, 8, 21, -3, -9, -4, 11, -7, 4, -8, -9, 2, 2, 10, 1, -15, -12, -2, 1, 11, 3, 12, 2, -7, 18, -14, -13, 2, 14, 11, 12, -17, -3, -7, 3, 2, -14, -11, 20, 8, 8, -11, -1, -10, 14, -4, 1, -8, 3, 2, 0, -2, 7, 1, 9, -13, 1, -10, -14, -4, -4, -11, 9, -12, -24, -2, 10, 1, 6, -5, -23, -6, -7, 1, -2, 0, -3, -7, -7, -24, -8, 10, 2, 0, -14, -5, -1, -11, 10, 8, -11, -5, -7, 4, -27, -8, -6, 2, -1, -13, -5, -16, -2, 2, 3, 14, -9, -19, -22, -10, -10, 2, -33, 7, 22, 18, -1, 11, -6, -2, 6, 11, -1, -3, -20, -15, 3, 12, 14, -6, 14, 9, -5, -14, -22, 1, 4, 22, -3, -10, -19, -22, -17, -12, -26, 11, 8, 10, 2, 17, -27, -4, -6, 8, 2, -1, -10, 4, 6, 1, 0, -5, 10, 9, 10, -2, -7, -3, 2, 20, -7, -5, -19, 20, -3, -6, -5, 4, -3, -2, 4, 8, -11, -7, -7, 4, 2, -2, 10, -15, 11, -7, 14, -3, -3, -12, 19, -19, -18, -3, -4, 17, 6, -3, -3, -13, -7, 0, -15, 8, -1, 0, -6, -2, 0, -19, -13, -6, 17, 8, -15, -8, 0, -15, -3, 3, -1, -5, 11, -3, -13, 5, -2, 2, -19, -6, -8, -6, -11, 19, 2, 6, 15, -2, -4, -6, -5, -7, 12, -8, 8, -2, 10, -6, 12, -10, -10, 8, 10, 2, 43, -2, 8, 8, -6, 2, -2, 8, 2, 3, -5, 15, 13, 8, 13, -16, -2, -3, 20, -2, 1),
    (7, -16, -9, 8, 2, 1, -9, 15, 5, 0, -10, -2, -5, -32, 5, 9, 3, 4, 9, 7, 9, 6, -6, -7, -3, 8, -26, -28, 10, 6, 2, -14, 5, -9, -12, 2, 2, 20, 0, -5, -15, 3, -18, -6, -12, -24, -12, 14, 10, -11, -2, 11, 12, 13, -5, -7, -7, 1, -1, -7, 1, 0, 4, -17, -9, 2, 4, 1, 9, -9, 6, -2, -30, 10, -14, -13, 2, -8, -28, 13, -20, -6, 8, 5, 11, 5, -5, -1, -20, 3, -5, 3, -22, -12, 1, -18, 5, -8, -3, -3, -15, 12, -8, -4, -22, -6, 6, 9, -10, 6, -2, 5, 3, -14, 7, 11, 7, -1, 13, 2, 10, -5, 2, -13, -19, -20, -4, 2, 1, -2, -5, -8, -1, 13, -12, -6, -8, -18, 17, 21, -14, 2, -14, 1, -2, -2, 15, 11, 18, 1, 15, 0, 5, -10, 1, 6, -17, -15, 1, 22, -2, 10, -2, -8, -2, 9, -6, -1, -2, -3, 11, 13, -2, 7, -4, -14, -1, 4, 7, 0, 2, -8, 5, 7, -9, -2, 6, 15, 6, -11, 4, 8, 3, -4, 1, -16, 7, -7, -10, -12, 4, 3, 2, 9, -16, 4, 1, -10, 5, 1, -1, -6, -19, -1, 7, 1, 11, -6, 8, 8, 3, 5, 3, 7, 7, -5, -2, -3, 5, -2, 2, 6, 12, -6, 8, 12, -8, 4, -1, -8, -4, 6, 3, -15, -4, 9, 0, -2, -3, -7, -8, 3, 22, -1, 10, 3, 1, -6, 3, -2, -2, -3, -32, -5, 6, -3, -13, 12, -11, -17, -6, 0, -4, -28, 1, -10, -12, -4, 3, -14, -11, 0, -15, 9, 18, -7, 7, -1, -6),
    (14, -5, 1, -14, -6, -5, 8, 5, 1, -5, -6, 0, 3, -2, 6, -6, -14, 22, 1, -15, -14, -14, -15, 10, -7, 4, -6, 2, -9, 2, -3, 22, 11, -2, 6, -8, -9, -17, 2, 2, 8, 11, 0, 6, 22, 0, 10, -10, -19, 5, -9, 3, -7, -16, -18, 13, -6, 2, 13, 2, 11, 9, -1, 19, 7, 4, -2, 2, -2, 0, 0, 6, -9, 8, 14, 0, 12, -6, 14, 2, -13, -2, -3, 6, -2, -12, -3, 5, -2, -10, 8, -6, 7, 4, -2, -1, 7, -12, -16, -11, 12, 3, 10, -4, 10, 9, 2, 5, -2, -7, -16, 10, -9, 5, -10, -17, -4, -21, -6, -10, -15, -2, -23, -14, -10, 12, 8, -8, 10, -2, -1, 3, 11, 6, 14, -4, 17, 14, 4, -6, 15, -7, 2, 5, -8, 6, -12, -27, -8, -2, -14, 15, -14, -2, 8, 10, 30, 14, 0, 5, 18, -3, 4, 17, 0, -4, 7, 4, 16, 18, -2, -11, 0, -7, 14, 18, 4, -15, -8, 1, -16, -5, -16, 4, -6, -7, 6, -1, 26, 17, 9, -9, -17, 12, -28, 3, -19, 6, -10, -8, 3, 1, -20, 3, -14, -21, -6, 9, -15, -5, -13, -19, -24, -4, -7, -28, -25, -7, -3, -28, -4, 9, 12, -2, 9, 6, -8, 5, 0, 7, 14, -11, 12, -3, 1, 7, 3, -13, 2, 4, 6, 2, 12, 11, -21, -2, -1, -18, -6, 6, 10, -1, 10, 7, 11, 6, -16, -9, -2, -4, -2, -3, 17, -5, 5, -15, -13, 4, -7, -8, 1, 2, -5, 11, -3, -1, -22, -2, -18, -12, -17, -5, -17, -5, 7, -5, -14, -8, -12)
  );
  ----------------
  CONSTANT Flatten_1_Columns : NATURAL := 2;
  CONSTANT Flatten_1_Rows    : NATURAL := 2;
  CONSTANT Flatten_1_Values  : NATURAL := 32;
  ----------------
  CONSTANT NN_Layer_1_Activation : Activation_T := relu;
  CONSTANT NN_Layer_1_Inputs     : NATURAL := 128;
  CONSTANT NN_Layer_1_Outputs    : NATURAL := 10;
  CONSTANT NN_Layer_1_Out_Offset : INTEGER := 6;
  CONSTANT NN_Layer_1_Offset     : INTEGER := 0;
  CONSTANT NN_Layer_1 : CNN_Weights_T(0 to NN_Layer_1_Outputs-1, 0 to NN_Layer_1_Inputs) :=
  (
    (8, 28, -47, -3, 7, 20, -29, 20, 13, 11, -69, -52, 27, -23, -38, 24, 4, -11, 27, 4, -21, 14, 47, -1, 10, -27, 21, -27, -20, 39, -93, 34, 14, 5, 24, 7, -23, 21, 14, 24, -8, -43, -56, -32, 3, 3, -2, 20, 20, -37, 51, 2, -22, 4, 35, 34, -21, 3, 9, -12, 12, -11, -65, -27, -14, 33, -43, -21, 5, -42, -17, 38, -17, 85, -30, -29, 31, 19, 13, 29, -20, -12, -17, -12, -30, -5, 10, -52, 5, 4, 32, -18, -11, -10, -24, -5, 8, 12, 7, 2, -15, 12, -16, -7, 24, -8, -13, -10, -7, -10, -19, -2, -11, -18, 7, -14, 9, 12, -18, -61, -23, 24, 12, -29, -12, 1, -26, 5, 20),
    (-92, -12, 1, -2, 12, -41, -33, 37, 18, 31, -30, -31, 19, 36, -2, -41, 19, -12, -27, -3, -8, 12, -9, -35, -45, 6, -73, 29, 52, -19, 3, -12, -41, -36, 5, -9, 7, 8, -20, 33, 4, 19, -46, -8, 20, -59, -17, -6, -14, -7, -27, -31, -20, 17, 9, -7, 2, -11, 13, 21, 17, -12, -16, -19, 6, 3, 17, -12, -7, -2, 20, -6, -5, 2, 10, 3, 22, 0, 5, -6, -6, -4, 20, -12, 26, -13, 19, 12, -10, 3, -9, 16, 24, 5, 32, 4, 13, 13, -9, 16, -2, 12, -1, -5, 9, -3, -7, -17, 10, -11, -10, -1, 0, -3, -17, 0, 4, 9, 31, 17, -12, 25, -3, 4, -3, 26, -17, -4, 22),
    (-3, 8, -13, 12, -8, -24, -60, -43, -3, 6, -9, 35, 14, 13, -44, -44, -6, 0, 23, -23, -19, 4, -24, -29, -22, 28, -22, -12, 20, 20, -27, 30, 3, 4, -10, 12, 0, -39, 11, -22, 3, -4, 1, 35, 12, 2, -11, -39, 0, -12, 15, 20, -40, -29, -32, -46, 1, 18, -3, 18, -17, 6, -20, -8, -5, -3, 3, 18, -29, 27, 0, -9, 31, 7, 1, 5, -13, 16, 6, -15, 6, 11, 35, 3, 4, 11, 1, -17, 10, 16, -25, 24, 17, 9, -5, 17, 5, 18, -10, -19, 6, 8, -19, 9, 0, 30, 4, 3, 4, 11, 5, -12, -10, 22, 8, 19, -48, 9, -8, 31, 30, -20, -15, 18, 20, 15, 12, 9, 36),
    (12, 22, -47, -24, -20, -28, 32, 19, 6, 8, 44, 5, -19, -30, 34, -12, -28, -28, 26, -44, 37, -12, -41, -4, 27, -19, 18, 25, -18, -16, 28, -23, 27, 18, 33, -11, -4, 27, 20, 24, 9, -27, -16, -10, -15, -17, 18, 11, 3, -19, 48, 0, 12, -16, 29, -7, -1, 19, 20, 3, -16, 14, -3, 11, -19, 12, 5, -63, -4, -17, -3, -22, -20, 4, 28, -4, -16, -11, 21, 1, -36, -20, -35, -28, 20, -4, -16, 36, -15, -29, 47, -24, -23, 20, 56, 33, 12, 1, 8, 22, 5, 4, -2, -19, -2, -7, 3, -15, -19, -3, 2, -13, 29, 7, -29, -12, 14, -12, -16, 31, -18, 2, 34, -10, -27, 0, 3, 15, -22),
    (5, -32, 12, 36, -36, 52, -15, -38, -5, -60, -21, 3, -48, -29, -42, 33, -20, 2, -4, 20, -3, -51, -5, 28, -24, 24, -21, -37, -19, -16, 13, 18, -18, -34, 11, 36, -9, 18, -22, 4, 5, -35, 2, 9, -2, 44, -15, 25, 32, 5, -15, 11, -8, 0, -14, 19, 31, 8, -3, -12, -22, 33, 28, -35, -25, -14, -1, 2, -14, 13, 1, -2, 20, -2, -12, 12, -12, -21, -16, 8, 15, 4, 4, -8, -14, 17, -8, 18, 12, 5, -17, 20, 3, 8, -16, 1, 0, 15, -1, -8, -1, 1, -43, 33, 3, 21, -14, 9, -5, 8, 21, -8, -14, 6, -26, 3, -12, 14, 6, -6, 13, -18, -7, 5, 9, 11, 27, -27, 49),
    (-39, -21, 8, 36, 30, 36, -13, 18, -54, -74, -8, -69, -4, -26, -19, 28, -44, -28, 17, 13, 37, -53, -28, -19, 11, -19, 22, 1, -12, -3, 18, -44, -45, -19, 21, 36, 1, 3, -31, 14, -21, -33, 7, 12, -11, 18, 26, 17, 17, 3, -24, -22, 5, -34, -57, 13, 4, -18, 7, 14, -21, -6, 29, -38, -8, -18, 4, 5, -43, 13, 5, -39, -23, 30, -47, -3, 22, -19, -40, -28, 18, 3, 35, 14, 27, 6, 27, -12, 4, 14, 21, 12, -22, -3, 20, -54, 25, 19, -19, -10, -13, 12, -17, -15, -15, -28, -10, 20, 3, -28, -11, -19, -5, 10, 4, 7, 18, -39, 14, -7, -7, -11, -14, -11, 9, 9, 28, -33, -100),
    (4, 28, -21, -54, -50, -20, -7, -31, 44, 28, 4, -2, -12, 35, 20, -55, 29, -14, -34, 5, -53, 33, 28, 36, 4, 12, -16, -27, 28, 12, -6, 24, 22, -3, 35, -20, -43, -2, -3, -12, -4, -3, 3, -21, -13, -33, 30, -30, 24, -2, 7, 14, -13, 16, 27, 36, 0, 5, -6, -13, 4, -3, -30, 37, -14, 23, 17, -59, 20, -24, -10, 31, -4, -26, 27, -24, -7, 28, 16, 10, -27, -20, -56, -18, -32, -19, 18, -9, 2, -10, 31, -41, -4, 5, 50, 32, -1, -13, 16, 19, 0, -5, -2, 12, 11, -35, 0, -20, -19, -11, -12, -10, 14, -18, -31, -30, -3, -37, 16, 15, -13, 5, 1, -25, -9, -6, -24, 4, -76),
    (11, 38, 20, 12, -2, -27, 3, -28, -5, -3, -35, -5, 30, 2, -34, -20, 12, 22, 4, 12, 20, 29, 4, -19, -19, -30, -4, -26, -19, -28, 4, -4, 26, -1, 11, 20, 9, -31, 7, -1, 5, -11, -29, 16, 14, 14, -3, 3, 4, 17, -5, 15, -2, -14, -20, -5, 4, -24, 5, -21, -11, 4, -4, -16, 5, -3, -3, 20, -18, 11, 15, -17, -19, -27, 2, 4, 19, 4, -28, -12, 19, 13, 5, 4, 27, 0, -13, -10, 16, 15, 16, 18, -28, 10, -26, -4, 21, 7, -7, -5, 5, -4, -17, -24, -14, 39, -12, 10, 1, 13, 9, -17, 1, 17, -5, 11, 17, 6, -13, -14, 8, -7, 14, 6, 4, 13, -1, -17, 39),
    (28, -21, 21, -28, -36, -11, 29, -27, 5, 13, 31, 29, -44, 12, 4, -34, -34, 28, -18, -5, -12, 3, -33, -13, 28, -3, 29, 12, -28, -20, 28, 3, 20, 11, -10, -12, -30, -17, 4, 5, 2, 13, 26, 12, -23, -3, 15, -48, 11, 38, 11, 11, -36, -10, 27, -35, 5, 4, -3, 13, -7, -8, 13, 4, -36, 12, 25, -57, 14, -19, -3, 35, 12, -34, 28, -33, -30, 28, 36, 10, -15, 3, -22, -14, 3, 0, -21, 12, -2, -22, -5, -27, -11, 10, 42, 29, 11, -11, 4, 6, -1, 6, -13, -1, 9, -21, 10, -7, -15, -13, 8, -8, 14, 10, -22, -16, -13, -20, -33, 26, -7, 13, 5, -10, -16, 5, 27, 4, -29),
    (-12, -36, 12, 34, 29, -16, -34, 12, -60, 28, -3, 5, -20, 35, -18, -31, -25, 4, -24, 37, 4, -36, 27, 52, 41, -31, -4, -5, 20, -34, -12, -67, -22, -18, -14, 23, 2, -31, -4, -8, -25, 27, 22, 14, -17, -14, -4, -19, 7, -2, -64, 24, 8, -19, -30, 6, 21, -3, -17, -12, 21, 12, 3, 0, -3, -36, -9, 16, -13, 4, 20, -18, 16, 29, -19, 3, 4, -10, -33, -27, 29, -27, 22, 12, -22, -15, 32, -52, 35, 7, -32, -1, -1, -35, -1, -57, -5, 14, -15, -21, -52, -1, -2, 5, 13, 8, -28, 11, 13, -22, 6, 4, -25, 8, -1, 4, -29, -18, 4, -25, 8, -15, -46, 1, 29, -22, 3, -37, 10)
  );
  ----------------
END PACKAGE CNN_Data_Package;
