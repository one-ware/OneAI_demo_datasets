library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.numeric_std.all;
use work.CNN_Config_Package.all;

PACKAGE CNN_Data_Package is
  CONSTANT Layer_1_Columns    : NATURAL := 128;
  CONSTANT Layer_1_Rows       : NATURAL := 128;
  CONSTANT Layer_1_Strides    : NATURAL := 1;
  CONSTANT Layer_1_Activation : Activation_T := relu;
  CONSTANT Layer_1_Padding    : Padding_T := same;
  CONSTANT Layer_1_Values     : NATURAL := 1;
  CONSTANT Layer_1_Filter_X   : NATURAL := 3;
  CONSTANT Layer_1_Filter_Y   : NATURAL := 3;
  CONSTANT Layer_1_Filters    : NATURAL := 8;
  CONSTANT Layer_1_Inputs     : NATURAL := 10;
  CONSTANT Layer_1_Out_Offset : INTEGER := 3;
  CONSTANT Layer_1_Offset     : INTEGER := 1;
  CONSTANT Layer_1 : CNN_Weights_T(0 to Layer_1_Filters-1, 0 to Layer_1_Inputs-1) :=
  (
    (-24, 8, -66, 45, -22, 46, -5, -8, -55, 0),
    (-15, 26, 5, 15, 44, 7, 19, 70, 8, 2),
    (14, 63, 18, 29, -16, 6, -35, -43, -53, 4),
    (49, 48, 19, -20, -11, -5, 4, 0, 49, -5),
    (16, 1, 9, 57, -50, 25, 0, 13, 15, -6),
    (31, -1, -26, 47, 35, -30, 27, -16, -32, -7),
    (37, 75, -1, 18, -34, 12, 26, 38, -46, -9),
    (10, -28, -34, -8, 6, 78, 11, -25, 45, 0)
  );
  ----------------
  CONSTANT Pooling_1_Columns      : NATURAL := 128;
  CONSTANT Pooling_1_Rows         : NATURAL := 128;
  CONSTANT Pooling_1_Values       : NATURAL := 8;
  CONSTANT Pooling_1_Filter_X     : NATURAL := 2;
  CONSTANT Pooling_1_Filter_Y     : NATURAL := 2;
  CONSTANT Pooling_1_Strides      : NATURAL := 2;
  CONSTANT Pooling_1_Padding      : Padding_T := valid;
  ----------------
  CONSTANT Layer_2_Columns    : NATURAL := 64;
  CONSTANT Layer_2_Rows       : NATURAL := 64;
  CONSTANT Layer_2_Strides    : NATURAL := 2;
  CONSTANT Layer_2_Activation : Activation_T := relu;
  CONSTANT Layer_2_Padding    : Padding_T := same;
  CONSTANT Layer_2_Values     : NATURAL := 8;
  CONSTANT Layer_2_Filter_X   : NATURAL := 3;
  CONSTANT Layer_2_Filter_Y   : NATURAL := 3;
  CONSTANT Layer_2_Filters    : NATURAL := 12;
  CONSTANT Layer_2_Inputs     : NATURAL := 73;
  CONSTANT Layer_2_Out_Offset : INTEGER := 4;
  CONSTANT Layer_2_Offset     : INTEGER := 0;
  CONSTANT Layer_2 : CNN_Weights_T(0 to Layer_2_Filters-1, 0 to Layer_2_Inputs-1) :=
  (
    (29, 8, 20, -12, -17, 59, 25, -22, 29, 32, 24, -20, -41, 53, 18, 3, 4, 9, 8, 7, 6, 7, 11, 4, 46, -4, 13, -9, 3, 37, 1, -9, 35, 37, 22, -32, -21, 63, 1, 1, 9, 28, 29, 1, 10, 18, 7, 0, 20, 9, 21, 3, -45, 46, 8, -10, 43, 11, 20, 10, -39, 28, 20, -5, 4, 18, 25, -36, 6, -6, 24, -6, -10),
    (7, 49, 44, 8, -2, 35, 36, 12, -18, 18, 2, 9, -9, 35, 29, -35, -21, -36, -7, -26, 7, 4, -22, -13, -15, -5, 41, -23, 11, 65, 41, -3, -5, -7, -12, -22, -25, 18, 11, -31, -27, -29, -35, 12, -16, -51, -28, 6, 2, -34, 38, -1, -4, 9, -28, -6, -66, -36, -12, -22, 12, -38, -57, -4, -59, 37, -48, 47, 7, -47, -7, 39, 1),
    (65, 21, -25, -34, -17, 4, 6, 2, 25, 25, -11, -18, -9, 40, -5, 30, 13, -5, -54, -2, 12, -16, -34, -27, 70, 71, -13, 28, 28, 6, -21, 18, 68, 53, 18, 10, -10, 12, 1, 34, 33, 36, -12, 36, 4, 12, -8, 29, 54, -21, 0, -6, -20, 12, -3, -5, 56, 11, 20, -25, 10, 9, 10, -19, 21, 4, 20, 22, 23, -9, -7, -14, -9),
    (-31, 21, -90, 12, -10, -20, -31, -16, -60, -8, -69, -22, 19, -27, -15, -16, -16, 19, -29, 2, -19, -6, -28, -29, 40, 36, -5, 42, 37, 11, 10, 11, 16, 31, -20, 9, 0, -5, -13, 12, 22, -17, -50, 22, 11, -6, -27, 12, 8, -6, 33, 15, 3, -22, -29, -15, 6, 4, 14, 36, 5, -18, -12, -11, 1, 37, 14, 56, 44, -27, -3, 12, 3),
    (49, -14, -9, -20, 11, -8, 9, 5, -23, -45, 19, -14, 4, -42, -52, -43, -45, 10, 37, 24, 46, -47, -3, 23, 39, 25, -18, 9, 53, 25, 33, 27, 19, -27, -57, -7, 3, 2, -6, -68, -39, -30, 16, 26, -15, -31, -10, 8, 34, 48, -1, 33, 59, 30, -4, 57, 12, 5, -36, -38, -18, 10, 18, -33, 8, -23, -27, -28, -27, 18, -8, -1, 15),
    (-29, -35, -21, -11, 21, -33, -37, -27, 18, 12, -69, 24, 0, -42, -36, -11, 50, 12, -30, 47, 18, -16, 20, 15, -38, -4, -50, -8, -31, -34, 4, -40, 33, 4, -87, 28, 17, -19, 6, -4, 93, 5, -34, -9, 45, 13, 10, 46, -36, -4, -50, -14, -32, -33, -31, -8, 11, -10, -53, -3, 22, -12, 23, 14, 36, 23, -25, -1, 38, 31, 43, 24, 4),
    (24, 6, -34, 7, 33, 7, 40, 13, 23, 36, -60, 31, 21, 6, -5, -6, 25, -13, -49, 15, 6, -4, -1, 6, 57, 5, -41, 23, 22, 18, 11, 4, 44, 3, -70, 27, 15, -4, 24, 8, 46, -2, -85, 11, 13, -23, -23, -5, 49, -19, -47, 12, 10, 4, 9, -13, 26, 5, -46, 32, 10, -10, 13, 4, 46, -13, -48, 47, 21, -12, -30, 22, 5),
    (-5, -28, -54, -29, -17, -57, -8, -17, 42, 40, 32, 7, 48, 47, 3, 26, 9, -23, -16, -24, -7, 21, 8, -46, 1, 4, -54, 1, -36, -43, -23, 20, 56, -7, 33, 28, 20, 44, 1, 50, 15, -28, -16, -6, -34, -15, 16, -78, 11, -10, -45, 4, -28, -9, -43, 28, 31, 4, 8, 22, -4, 25, 20, 21, 4, -50, -9, 13, -4, -16, -8, -22, 4),
    (23, 19, 15, 52, 55, 18, -4, 10, 32, 45, 20, 51, 0, 7, 6, 34, -5, 48, -13, 23, 4, -6, 28, 46, 3, -46, 15, 0, -3, -2, 7, -7, -2, -7, 44, 13, 14, 1, -26, -1, -36, 5, 36, 10, 10, -3, 8, 9, -70, -39, 14, -6, -4, -8, -12, -23, -98, -34, 37, -9, -45, 3, -45, -44, -68, -39, 28, -32, -12, -4, -9, -13, 5),
    (28, 14, -21, 25, 29, -7, 21, 2, -23, -16, -21, 38, 23, -8, 29, -25, -22, -25, -31, 22, 5, -2, 38, -43, 38, -13, -29, 34, 28, -15, 16, 0, 6, -15, -38, 26, 30, -29, 36, -30, -12, -39, -33, 37, 29, -13, 36, -51, 29, -5, -27, 33, 35, -15, 25, 4, 20, -18, -26, 17, 2, -22, 26, -9, 14, -45, 0, -8, -11, 8, 5, -33, 2),
    (3, 0, -11, 2, 12, 27, 32, 18, -3, 41, -12, -32, -5, 11, -2, -15, -6, 35, -43, 12, 24, 27, -1, 18, -38, 17, -2, -4, -17, 0, 35, 1, 7, 3, -8, -6, 4, 0, -3, -21, -40, -4, 13, 2, 38, -26, 12, 2, 2, 52, -29, 0, 47, -12, 2, 21, 19, 46, -21, 15, -7, -28, 11, -10, -12, 37, -29, 27, 21, -19, 6, 27, -6),
    (-15, -8, 10, -13, -23, -46, -16, -41, 45, -2, -27, -1, -18, 7, -34, -10, 21, 34, -8, -2, 16, -3, -24, -41, 15, 0, -13, -24, -11, -38, -40, -50, 34, -25, -9, -32, -18, 11, 24, 12, 3, 38, -37, -11, -25, 3, -1, 8, -22, 20, 44, 16, -14, 23, 4, -46, 17, -11, -9, 41, 8, -26, -45, 28, 13, 1, -45, 25, -16, -2, -10, -37, 1)
  );
  ----------------
  CONSTANT Layer_3_Columns    : NATURAL := 32;
  CONSTANT Layer_3_Rows       : NATURAL := 32;
  CONSTANT Layer_3_Strides    : NATURAL := 2;
  CONSTANT Layer_3_Activation : Activation_T := relu;
  CONSTANT Layer_3_Padding    : Padding_T := same;
  CONSTANT Layer_3_Values     : NATURAL := 12;
  CONSTANT Layer_3_Filter_X   : NATURAL := 3;
  CONSTANT Layer_3_Filter_Y   : NATURAL := 3;
  CONSTANT Layer_3_Filters    : NATURAL := 16;
  CONSTANT Layer_3_Inputs     : NATURAL := 109;
  CONSTANT Layer_3_Out_Offset : INTEGER := 6;
  CONSTANT Layer_3_Offset     : INTEGER := 0;
  CONSTANT Layer_3 : CNN_Weights_T(0 to Layer_3_Filters-1, 0 to Layer_3_Inputs-1) :=
  (
    (-23, -7, 20, 0, 22, 5, 23, 28, -4, 4, 17, 21, 12, 16, 8, -11, 24, 1, 12, 10, -26, -4, 4, 50, -5, 14, -12, 0, -11, -3, 5, -27, -25, -20, 12, 18, -3, -9, 20, 40, -5, 35, -1, -20, 5, 23, -4, -2, -26, -4, 61, 46, -16, 19, 27, -61, 37, -2, -20, -9, 35, 19, 50, 41, -22, 9, 5, -42, 22, 31, -21, -29, -39, -25, -55, -38, 49, -4, -36, 20, -20, -20, -29, 35, -27, -14, -49, -17, 28, -42, -33, -17, -1, -36, 35, -3, -1, 15, -26, -49, -12, -19, -34, -11, 2, -18, -17, 11, 4),
    (11, -40, -21, 25, -13, 4, -2, -1, -12, -5, -4, 13, 16, -45, 17, -16, 6, 21, 34, 19, -41, 41, 22, -4, 47, 16, 4, -29, 4, 39, 17, 23, -22, 21, 36, -36, -48, -50, -18, 4, -29, -13, -32, -39, -5, -16, -3, 12, -20, -80, 6, -14, 36, 2, 39, 26, -21, -1, 2, 12, 28, -38, 12, 30, 48, 28, 21, 19, -16, 10, 16, 41, -9, -31, -31, -23, -36, -20, -42, -15, -10, -7, -33, -34, -15, -70, -23, 16, 7, -11, 12, 9, -2, -8, -13, 19, -12, -15, 23, 20, 62, 29, 30, -16, 4, -1, 12, -10, 1),
    (20, -40, -3, 19, 34, 11, 3, -21, 6, -10, 8, -15, -26, 12, 19, 14, -38, 32, -13, -28, 0, 25, 3, -13, 8, 24, 31, -1, -44, 25, -17, -24, 6, 38, 23, -5, -11, -53, 18, 14, 30, -46, -23, -29, 26, -38, -16, 4, 5, -11, 19, 24, -3, -60, -36, -34, 44, -27, -21, -32, -7, 20, -45, -9, -54, -47, -52, -23, -12, -2, 0, 36, 1, -28, -3, 35, 11, 8, -14, -24, -13, -73, -16, -13, 5, -16, 11, 2, -26, -15, -20, -63, -5, -26, 12, 29, -6, 19, 10, 1, -34, -5, 12, -15, -19, -40, 15, 36, 4),
    (37, 37, 18, 31, -14, 19, 19, -2, 10, 28, -8, -20, 15, 46, 31, -3, -78, 2, -4, -7, 26, 15, 12, -51, 9, 33, -37, -28, -92, -16, -21, 6, 10, 18, 6, -8, -3, 6, -38, -12, -50, -45, -45, -45, -2, 9, -4, 8, -23, 12, -49, -1, -82, 3, -25, -34, -6, -25, -28, 21, -28, 45, -14, -4, -37, 19, -4, 9, -39, -34, 10, 14, -33, -17, -36, 9, -79, 3, -6, -21, 20, -31, 11, 31, -1, 26, 16, -17, -54, 11, 28, -25, -33, -12, -11, 41, 30, 22, -12, 11, 8, 21, 12, -7, -9, 29, 38, 24, 6),
    (-12, 6, -8, 8, 6, 0, -29, -15, -51, -73, -1, 9, -38, -55, -38, -21, 33, -24, -10, 2, -12, -61, -21, 30, 2, -33, 1, -31, 30, -13, -14, -15, 4, -14, -4, -2, 4, -12, 12, 22, -11, -7, 42, -45, -8, 13, 7, 15, -11, -45, 4, 19, 7, -12, 40, -20, 17, 12, 13, 22, -37, -38, 20, 49, 20, -5, 25, -19, -38, 14, -17, 4, 17, -1, -4, -2, -7, -5, 0, 2, -12, 20, 20, 7, 3, -38, -5, -4, 8, -11, 29, -27, -5, 0, 26, -10, 1, -34, 11, 37, 23, -7, 22, 1, 28, -14, -1, 2, 1),
    (-27, 37, 9, -11, -15, 28, 25, 46, -6, -3, 3, -13, -25, 53, 20, 5, -28, 33, -6, 57, -12, 44, 29, 25, -26, 22, 19, 8, -13, 5, 0, 12, 2, 31, 42, 48, 3, 60, 20, 10, -36, 29, 6, 11, -12, 41, 10, 3, -20, 72, -8, -4, -52, 29, -3, 48, -12, 52, -2, 37, -19, 18, -13, -36, -15, 4, 11, 31, -20, 38, -20, 31, -14, 40, -17, 12, -11, 5, 0, -24, -4, 28, -3, -40, -12, 28, -26, 5, -36, 1, -8, -16, -13, 23, -12, -8, 11, 3, -11, -13, -3, 20, -9, -26, -15, 11, -16, 11, 1),
    (-15, -38, -25, -45, 10, 5, -24, -6, 26, -25, -21, 5, 11, -43, 5, 16, -6, -4, -1, -20, 5, 0, -20, -3, 10, -9, 14, 25, -36, -4, -7, -44, 11, 32, -8, -1, 9, -35, -17, -6, 25, -16, -23, -23, -14, 9, -12, -15, -28, -66, -43, -20, 26, -19, -30, -42, -5, -25, -10, -1, -3, -23, -17, -49, 13, -22, -15, 18, -9, -7, -4, 21, 20, -49, -1, -9, 21, 4, 51, -31, 13, 32, 27, 2, 5, -51, 8, 15, 33, -4, 47, -38, 30, 15, 19, 22, 10, -23, -20, 35, 19, 11, 19, -3, 12, 8, 20, 1, 13),
    (-18, 15, 10, -30, 3, -13, -20, 6, -2, -36, 15, -18, 12, 12, 3, -33, 11, -5, -17, -20, 6, -20, 17, 10, -6, -10, 13, 8, -3, 13, -13, 0, -3, -12, 28, -7, 14, 6, 13, -29, -4, -7, -5, -14, -20, -32, 16, -2, 17, 32, 4, -18, -18, -8, 8, -13, 16, -21, 11, -8, 35, 18, -3, 30, -7, 32, 19, -2, 4, -27, 59, -12, 2, 23, 15, 11, -42, -1, 13, 13, -12, -31, 4, -25, 31, 20, 4, -13, -25, -4, 29, -33, 5, -17, 11, 26, 27, 5, -3, 24, -14, 30, 46, -49, 15, -18, 36, -28, -10),
    (-13, 12, -41, -30, -2, -13, -25, -29, 4, 13, -9, 2, -4, -18, -27, -12, -10, -33, 9, -70, 15, 26, 20, -20, 14, -30, -5, 19, 12, -19, 54, -42, 42, 9, 7, 14, 5, -8, -19, -21, -28, 8, 4, 0, -23, 15, -26, 51, -15, 2, -37, -11, -3, -30, 16, -38, 8, 34, -23, 17, 3, -2, -32, -19, 13, -5, -3, -23, -2, 22, 20, -16, -1, 0, -18, 21, -27, 15, 16, 11, -17, -31, -16, -7, 17, 5, -3, -15, -37, 17, 5, 10, -39, -23, -9, -7, -27, 4, -2, -3, -33, 0, -34, 39, -44, 37, 22, 29, 2),
    (-16, -2, -15, -15, 27, -7, 17, -12, 5, 16, -21, -29, -15, 3, -19, 8, 13, 2, -18, -19, -43, 2, -4, -7, -13, 3, 3, 27, -6, 14, 14, -20, -42, 9, -13, 20, -25, 15, -41, 4, -2, 10, 2, 25, -38, -4, -1, 8, -9, 37, -8, 11, 3, 44, 29, 37, -66, 31, -20, 45, -11, 36, -4, -9, -10, 46, 40, 7, -45, 13, 17, 25, -20, 27, 2, -8, 5, 3, 12, 45, -53, 0, 5, 26, -14, 34, -9, 20, 0, 59, 16, 48, -30, 10, 22, 9, 21, 29, -5, 28, 8, 53, 17, 28, -5, 4, -1, 42, 7),
    (20, -27, -7, 28, 36, -12, 31, -10, 6, 31, -13, 6, 0, -69, 25, -5, 49, -7, 2, -15, -35, 13, 4, 18, -35, -35, -20, -12, 19, -37, -25, -16, -19, -8, -21, 1, 1, -24, 18, -29, 44, 15, 25, 27, -22, 37, -12, -12, -10, -64, 12, 19, 58, 31, 21, 28, -57, 19, 9, 17, 7, -24, -42, -36, 20, -29, 12, 23, -56, 21, -33, -7, 21, -14, -23, -2, 35, 6, 17, 34, -23, 21, 21, -18, -1, -20, 5, 16, 25, 47, 22, 50, -50, 25, 32, 11, -10, 10, -21, -15, 12, -17, 17, 9, -44, 20, -28, -4, 8),
    (28, -27, -8, 25, 11, -28, 35, -52, 10, -2, 40, 33, -1, -24, 25, 8, 0, -30, 7, -46, 11, -21, 5, 1, -8, -1, 13, -6, -7, -30, 0, 13, 1, -30, 17, -30, 25, -28, -7, 19, 22, -45, 36, -47, 14, -9, 36, -17, 33, -61, 28, 15, 38, -62, 6, -65, 25, -37, 1, -29, 15, -30, 10, 15, 4, -34, 5, -38, 7, -19, 24, -22, 13, -5, -3, -28, 9, -13, 12, -5, -34, -14, -12, -21, 19, -12, 20, -5, 22, -33, 12, -35, -8, -15, 8, -37, 23, -15, 11, 13, 8, 1, 14, -2, 4, -1, 27, -55, -4),
    (31, 13, 31, -18, 29, 63, 27, 19, -2, 26, 6, 9, 8, 12, 17, -15, 2, -6, 4, 42, -27, 44, -18, -1, -5, -24, -46, -15, -13, -13, -25, 59, 3, -17, 10, 57, 24, -2, 7, 8, 53, 53, 9, 56, -6, 26, 10, 6, -26, 13, -6, -35, 3, -25, 16, 45, -31, 5, -6, -19, -9, 8, -24, -22, 3, 43, -13, 30, -37, -11, -19, 22, 1, -12, 11, 8, 15, 42, -8, 30, -23, 38, 0, -8, -20, 13, -4, -10, 4, 17, -3, -1, 10, 13, -8, 30, 12, 15, -7, 3, -27, 36, -31, 68, -38, -64, 3, -7, 1),
    (5, 3, -6, 13, -39, -14, -12, -63, 20, 13, 31, -6, 0, 12, -27, 33, -84, -29, -1, -49, 6, 9, 21, -4, 34, -12, -12, 10, -48, 1, 7, -69, 32, 7, -12, -5, 20, 17, 17, 2, -11, -8, -2, -43, 36, -8, 41, 5, 14, -5, -12, 23, -24, -1, 5, -50, 31, -8, 37, -5, 12, -19, -5, 19, -8, -22, 0, -17, 36, -12, 6, 16, 17, 16, -4, 13, 12, -9, -13, 11, 26, -17, 15, 1, 30, -2, -5, -13, 18, -8, -7, -4, 24, -19, -16, -28, -9, -20, 11, -4, 27, -33, -27, 31, 27, -4, -35, -22, 1),
    (21, 43, -6, -12, -20, 19, -13, 29, -26, 4, 23, -7, 23, 59, 11, -22, -38, 48, 1, 64, -44, -6, 17, 16, -2, 34, -3, -2, -24, 25, -18, 43, -6, -6, -2, 11, 35, 40, 11, 10, -32, 20, 32, 8, -7, -4, 10, 5, 45, 46, 10, -2, -44, 67, -8, 53, -31, -21, 12, 20, 11, 21, 13, -20, -8, 38, -24, 27, -18, -2, -15, -31, 31, 7, 23, 8, 2, 1, 16, -6, -17, 12, 33, 31, 33, -6, 7, -10, -12, 29, -3, 34, -32, -12, -7, 48, 10, -20, -5, -4, 16, 8, 4, 20, 4, -20, -14, 31, -8),
    (-12, 22, 2, 5, -28, 15, -14, -5, 32, 23, 11, 26, 17, -13, 39, 49, 13, 17, 36, -35, 46, 15, -11, -28, -3, -20, 42, 22, 31, 19, 26, -42, 20, 1, -6, -44, -20, 11, -39, -11, 25, 2, -20, 46, -45, 1, -5, 28, -20, 7, -52, -38, 23, -28, -37, -18, 21, -19, -22, -10, -20, -14, -3, -16, 12, -8, -17, 20, 35, -2, 15, 0, 6, -10, 20, 33, 12, -18, 12, -31, 7, 11, 14, -26, -31, 2, 18, 18, 1, 4, 8, -34, -51, 4, 22, -13, -25, 31, -30, -16, -9, -6, -32, 28, -14, 8, 13, 11, -6)
  );
  ----------------
  CONSTANT Layer_4_Columns    : NATURAL := 16;
  CONSTANT Layer_4_Rows       : NATURAL := 16;
  CONSTANT Layer_4_Strides    : NATURAL := 2;
  CONSTANT Layer_4_Activation : Activation_T := relu;
  CONSTANT Layer_4_Padding    : Padding_T := same;
  CONSTANT Layer_4_Values     : NATURAL := 16;
  CONSTANT Layer_4_Filter_X   : NATURAL := 3;
  CONSTANT Layer_4_Filter_Y   : NATURAL := 3;
  CONSTANT Layer_4_Filters    : NATURAL := 24;
  CONSTANT Layer_4_Inputs     : NATURAL := 145;
  CONSTANT Layer_4_Out_Offset : INTEGER := 6;
  CONSTANT Layer_4_Offset     : INTEGER := 0;
  CONSTANT Layer_4 : CNN_Weights_T(0 to Layer_4_Filters-1, 0 to Layer_4_Inputs-1) :=
  (
    (-51, -39, 4, -21, -13, -11, -18, -44, 21, 0, 33, -20, -29, -39, -12, -33, -12, -6, 31, -4, 18, -7, 9, 1, 9, 7, 4, 1, -30, -35, -34, -7, -7, 2, 14, 20, -2, 41, 19, 22, -6, 18, -12, -13, 16, -2, -20, -8, 6, 24, -12, -17, -14, -4, -8, 11, -12, 17, 28, -40, 3, -7, -26, -22, 36, 14, 53, 18, -5, -4, 4, -11, -5, 36, 9, -22, 12, -1, -21, 5, 6, 7, 31, 68, 3, 33, 20, -23, -3, 5, 17, -30, 11, -5, 6, -4, 36, 16, 13, 59, -15, 8, -22, -13, -22, 52, -30, 27, 1, 32, 19, 28, 20, 26, 11, 31, -25, 11, -19, 8, 1, 33, -29, -23, 10, 18, -1, 36, -1, 0, 11, 22, -16, 33, 11, -35, -13, 12, -13, -47, -10, 0, -22, -11, 2),
    (35, -40, 26, 31, 13, 13, 10, 20, -17, -23, -27, -31, -20, -6, 26, -6, 28, -32, 32, 2, -1, -6, 4, 21, -7, -21, -16, 9, -12, 6, 30, 12, 13, 4, 2, -20, -22, 6, -8, 13, 55, -22, -4, 4, 12, -20, 9, 25, 5, -15, 4, 22, 13, 12, 30, 0, -41, -34, -35, 30, -13, -1, 16, 15, 11, -22, 16, 1, 20, 12, 26, 7, 13, -28, -23, 25, -12, 26, 18, 28, 20, -12, 13, -13, 4, 11, 4, 41, -20, -17, -5, -24, -4, 10, 23, 12, 7, 13, 1, 1, -19, -7, -4, 14, -36, -10, -10, -36, -8, -17, 17, 1, -5, 11, 1, 20, -27, 3, -31, -4, -34, 19, -19, -1, 3, -9, 29, 2, -3, 5, 13, 20, -29, 12, -42, -8, -3, 21, -13, -10, 0, 11, 22, -7, -4),
    (-22, -5, -17, -31, 1, -35, -3, 8, -25, -10, -6, -5, -21, -15, -22, -36, -6, -4, -14, -51, -20, -27, -7, -5, -49, -10, 17, -11, -28, 0, -31, -37, -28, 1, -58, -27, -10, -9, -2, 1, -46, -5, 21, 2, -6, -35, 11, -7, -12, 38, -27, -60, -13, -12, -9, 12, -23, 1, 30, -19, 7, -32, -21, -4, -27, 44, -3, -44, -18, -3, -1, -9, -17, 20, 21, 4, 17, -31, -18, -17, -53, 38, -16, -20, -6, 5, 8, 4, -36, 4, 26, -15, 18, -27, 0, -33, -1, 32, -29, -13, -13, -2, -11, 21, -15, 12, 37, -31, 33, 2, 4, 3, -23, 39, -26, -11, -4, 5, 0, -3, -20, 27, 43, -13, 30, -23, -6, -4, -23, 38, -47, 16, -9, 22, 4, 9, -5, 24, 32, -2, 11, -11, -8, -19, 7),
    (-20, 36, -28, 1, -14, 1, -9, 16, 16, 10, 0, 36, -12, 12, 2, -6, 4, 64, -22, -16, -9, -11, -25, 0, 21, 5, -27, 36, -13, 23, 5, 27, 19, 3, -13, -11, 11, -15, -8, -20, 24, -12, -29, 1, -13, 7, -12, 28, -19, 45, -38, -29, -2, -4, -20, 0, -6, 0, 36, 47, -6, 13, -22, -2, 10, 63, -25, -53, -13, -20, -23, 3, 22, -4, 27, 44, -7, 26, -32, 33, 15, 36, -4, -28, -12, -13, 1, -15, 27, -52, 14, 3, -12, -8, -13, 34, 4, 8, 6, -29, -12, -15, -15, -12, -10, -15, 28, 7, 21, 9, -5, 9, 0, -6, -4, -23, -21, -4, -16, 13, 5, -37, 48, 8, 24, 2, -1, 6, 4, -10, -4, 14, -8, 6, 3, 0, 3, -57, 12, -23, 4, -7, 19, 3, -4),
    (-13, -21, 0, 17, 7, -2, -14, 20, 7, 10, -10, -1, -15, -16, -8, -12, -27, 17, -22, -5, -27, 20, -42, -2, 19, 3, 21, -5, 11, 9, 28, -12, -4, 38, 3, 10, 2, 2, -16, 9, -11, 8, 13, 2, 4, 44, 34, 10, -52, 19, -22, 4, -59, 12, -30, 19, -10, 12, 4, -23, -4, -8, -8, -12, -20, 42, -47, -44, -96, -8, -48, -14, 10, 18, 24, -27, 29, -3, 34, 4, -5, 27, -15, -19, -20, 6, -19, 7, -6, 13, 17, -12, 14, 13, 40, 20, -17, 4, -22, -41, -84, -16, -44, -40, 25, -21, 14, -28, -25, -5, -14, -23, 4, 29, 3, -60, -52, -36, -21, -28, 26, -5, 6, -10, 8, -18, 7, 3, 9, 26, -4, -14, -5, -9, -9, 7, 5, 1, -13, -21, 8, -13, 28, 9, -5),
    (-24, -5, -8, 7, -16, 13, 4, 7, -61, 28, 13, -8, -9, -13, 21, -28, -32, -12, 9, 18, -16, 0, -10, 10, -29, 28, -12, -19, -3, -37, 37, -28, -26, -21, -4, -6, -10, -3, -7, -4, -66, 12, -18, -3, -1, -32, 0, -26, -5, 37, -28, 22, 20, 21, -56, 2, 29, 24, -15, 30, 9, 12, 20, 10, 28, 52, -16, 11, 27, 0, -19, 19, 17, 43, -31, 17, -19, 10, 6, 38, 25, 37, -4, 8, 17, -8, -10, 22, 14, 28, -37, 27, 3, 9, -5, 19, -22, 27, -20, -13, 17, -5, 10, -39, 14, -1, 17, -5, -11, 1, -33, 26, -11, -4, -19, -11, 36, 25, 29, -45, 13, 0, -18, -5, -1, -1, -27, 36, 3, -22, -19, -17, -5, 6, 7, -44, -6, -14, -37, -4, 5, -12, 1, 10, -1),
    (10, 12, 11, 0, 3, -14, 6, 27, -14, -5, 19, -8, -5, -17, -17, 3, -4, 29, 38, 21, -17, 4, 1, 32, 44, -4, 46, -4, 17, -6, 15, 7, -53, 16, -21, -36, -2, 8, -10, -13, 28, -1, 36, -12, 13, -8, -13, -33, 5, 1, 35, 35, -1, 21, -4, 25, -1, 13, 51, -34, 28, 3, 13, -28, -18, 19, 48, 24, -4, 28, -16, 11, 16, 20, 52, -26, 34, 5, 14, -52, -41, 34, -74, -20, -26, 20, -34, -37, 51, -3, 23, -3, 16, -15, 25, -51, -18, -21, 8, 28, 4, 2, 13, 12, 4, -9, 13, 7, 20, 9, 1, -5, -27, -8, 11, 12, -20, 22, -19, -3, 30, 13, 3, -11, 2, 16, 9, -29, -32, 16, -15, -8, -29, 12, -7, -3, 3, 12, -20, 5, -8, -9, 20, -18, 0),
    (21, 19, 2, -2, 11, -6, 6, 0, -20, 11, -21, 7, 15, -4, 8, 20, 30, -5, 7, -12, 1, -13, 12, -9, 25, -7, 3, 20, 5, 7, -18, 37, 10, -32, 17, -6, -17, -9, -9, -19, 27, -16, 28, -4, -5, -36, 12, 8, 52, -6, 35, 13, 32, -22, 30, -18, 2, -1, -12, 11, -26, 36, 12, 39, 41, -40, 39, -2, 19, -35, 27, -12, 45, 1, 4, 28, -23, -12, -5, 36, -3, -38, 21, 5, -4, -15, -16, -37, 24, -17, -13, 4, 6, -28, 13, -3, 13, -38, 19, -16, 11, -19, 18, 8, 4, -29, 13, 16, -12, 21, -2, 16, 9, -29, 7, -20, 5, -33, 5, -5, 34, -32, 23, -12, -15, 13, -18, 7, -28, -36, -7, -34, -26, -28, -17, -35, -13, -39, 41, -10, -4, -34, -21, -13, 4),
    (15, -10, 43, -21, -4, -58, 15, -37, 27, -10, -42, 20, -59, 3, -46, 8, -32, -15, -5, -8, 16, -17, 16, 2, 14, 12, -30, 5, -49, -22, -36, -13, 2, -29, 9, 9, 11, 34, -19, 0, 11, 25, -39, -9, -6, 12, 10, -12, -6, -13, 28, 45, 16, 41, 12, -4, -48, 29, -45, -40, -16, 7, -11, -38, -12, 1, 2, 67, -4, 52, -37, 5, -49, 48, -36, -9, 9, 23, 37, -39, 14, -12, 13, 21, -11, 20, -34, 3, -21, -4, -19, -7, -2, 18, 25, 4, -8, 4, -9, 31, -31, 18, -13, -2, -12, 28, -11, 4, 11, 25, 32, -1, 11, 24, 10, -19, -19, -18, -10, -4, -3, 15, -9, -4, 0, 23, 4, 19, 17, -23, 4, -30, -8, -21, 21, -4, 15, -35, -20, -5, 4, -32, -20, 19, -5),
    (-29, 4, -17, 13, 5, 29, -4, 11, -4, 3, -13, -11, 28, 2, 1, -7, -37, 23, -17, 15, -2, 61, -29, 20, -33, 25, 4, -18, 36, 31, 1, -21, -6, 39, -4, 10, -37, 40, -14, -6, -7, 8, 32, -17, 11, 16, 6, -5, -10, 6, 9, 20, -26, 28, -8, -12, -32, 32, -32, -19, 27, 1, 16, -26, -58, 39, -12, 1, -76, 38, -15, -13, -6, 36, -3, -5, 31, 5, 3, -33, -9, 30, -12, -21, -63, 4, -15, -33, -8, -12, 20, -3, 2, -29, -3, 2, 10, 4, 7, 5, -25, 7, 8, -13, 21, 28, -28, -5, 7, -15, 14, -7, 2, 11, -30, -31, -91, -2, -17, -22, 19, 2, -20, -3, 20, -4, -20, -10, 4, 25, 1, -24, -52, -34, -7, -15, -18, -22, -3, -20, 5, -20, -19, 5, 4),
    (-8, -4, -25, 20, -18, -4, -10, -8, 1, -9, 46, -13, -13, -20, 12, -12, -6, -4, -13, -14, -11, -24, -1, 2, -35, -20, -11, 9, 9, -12, 12, -13, 19, 8, 29, 2, -4, -46, -25, 13, -33, -13, -25, 18, -30, 30, 13, 13, -4, 11, -5, -8, -10, -18, 12, 5, -8, -21, 18, -34, -12, -14, -21, 4, 46, -3, 16, -38, -4, -32, 26, 14, -28, -54, 17, 20, -18, -12, -10, 12, 40, 7, 32, -5, -4, -4, 3, 37, -10, -38, 19, 38, -19, 4, 5, 28, 20, -11, 17, -26, 5, -32, 9, -17, 13, -18, -12, -27, -43, -31, -28, 10, 15, -12, 15, -20, 14, -21, 19, 5, -2, -36, -1, 11, -38, -4, -20, 22, 3, -13, 4, -2, 0, 20, 14, 33, 3, -13, 13, 12, 26, 12, 10, 8, 0),
    (11, -16, 27, -10, 4, -34, -17, -19, -28, -13, 7, -28, -41, 3, -34, -4, 27, -39, 21, 8, 14, -32, 21, -1, -11, -3, 23, 12, -34, -3, -39, 4, 31, -33, 22, 5, 12, 14, 17, 12, -19, 10, 3, -18, -10, 5, -21, 11, 19, -35, 22, -14, -38, -20, -44, -5, -15, -36, -24, 1, -48, -20, -48, -9, 22, -44, 37, 32, 27, 36, 4, 17, -21, -21, 0, 2, -7, 29, -34, 11, 16, -12, 23, 53, 48, 33, 18, 19, -13, 2, -4, 12, 7, 6, 14, 21, 15, -32, 25, 12, -10, 0, -11, -14, -11, -16, -51, -21, -29, 3, -4, -7, 14, -36, 24, 32, 9, 24, -2, 9, -12, -36, -46, -17, -5, 9, 20, 5, 4, -8, 23, 21, 8, 4, 4, 12, -19, 2, 2, -4, 4, 19, 5, 13, 0),
    (11, 21, 9, 22, -52, 4, 2, -2, 19, -5, -11, 5, -36, 18, 39, 3, 0, -15, 23, 25, -8, -4, 4, -18, 19, -6, -65, 1, -28, 25, 22, 3, -4, -55, 12, 4, -53, -6, -21, -37, 20, -26, -29, -32, -11, 9, 1, -7, -48, -42, 20, 16, 4, -31, 28, -18, 12, 19, -35, -12, -68, -28, -21, 15, -28, -52, 21, 9, 29, -30, 33, -4, 23, -18, -24, 6, -45, 10, -10, 1, -26, -54, 10, 12, 2, 3, 18, -25, -14, -49, 21, -25, -20, -22, -26, 0, -27, -20, -10, -1, 11, 2, 19, -4, -24, 20, -42, 13, -30, 29, 4, 7, 13, -60, 12, -1, 15, 4, 20, 8, -7, -24, -15, 14, -41, 0, -2, 33, 32, -35, -1, -42, 5, -5, 37, 13, -22, -21, 22, 8, -22, -16, 3, 10, 13),
    (16, 25, 12, 2, -4, -13, -39, -12, 24, -20, 3, 17, -11, 4, 12, 25, 17, 27, -4, -16, 12, -19, -11, 4, 79, -30, -4, 20, -29, 10, -10, 36, 16, 28, 3, 0, -3, -9, -29, 18, 77, -18, -16, 19, -4, 3, 4, 22, -28, -12, 19, -1, -5, 2, -9, -17, 18, -20, -24, -7, -48, -25, -39, 14, -50, -21, -41, -38, 26, 43, 26, -11, 39, -17, -21, 2, -4, 20, -17, 23, -32, -11, -43, -13, -18, 26, -12, -12, 36, 4, -18, 12, 4, 14, -9, 12, -11, 3, -12, 7, 10, 23, -16, -11, -1, 20, -24, -29, -12, 12, -6, -38, -15, 14, 6, 30, 11, 19, -42, -23, -30, 35, -30, -29, 27, 8, 13, -47, -4, -5, 5, 21, 3, 43, -42, -35, -3, 15, -7, -41, 23, -4, -11, -31, 1),
    (-26, 4, 0, 11, -3, 20, -10, -5, -7, 0, 30, -4, 30, 21, 3, -11, -21, 31, -11, 3, 1, 19, -3, -25, -3, 5, 45, -15, 22, -7, 27, -43, 20, -15, -15, -28, 41, -21, 30, 13, -40, -39, 1, -1, -11, -21, -35, -6, -28, -11, 6, 36, -45, 30, -17, 7, -18, 12, 27, -6, -2, -6, 28, -50, -52, 26, -26, -20, -51, 21, -28, -6, 46, -16, 26, -28, 4, 11, -6, -44, 19, -2, -11, -1, 28, -30, 3, -12, 25, -33, -29, 32, -32, 17, -34, 26, -20, -12, -11, 8, -62, 4, -70, 4, -14, 9, -14, -33, 4, -7, -3, -36, -31, 0, -33, -12, -63, -5, -21, -22, 4, -48, 4, -18, -11, -11, -9, -73, -16, -14, 11, -22, -33, 11, -4, -25, 1, -14, -17, -2, -20, 22, -27, 15, 18),
    (-6, 6, 5, 6, 11, 5, -6, 22, -12, 24, 9, 8, -4, 23, 23, 4, 3, 14, 0, 5, 11, 0, -24, 12, -3, 29, -22, 21, -24, 3, 28, -2, 9, 5, 9, 12, 11, -10, -18, 2, 0, 12, -47, 17, -19, 3, -5, 5, 29, 41, 2, -4, -5, -41, 19, -40, 13, 0, 13, -4, -19, 5, -32, 23, 12, 38, 6, 24, 15, -19, 15, -22, 34, -5, -31, 30, -55, -13, -7, 1, -11, -53, -3, 12, -2, 6, -28, -43, 21, -35, -29, -1, -51, 21, -7, 0, -52, 5, 0, -55, 3, -23, 16, -7, 12, -2, 32, -4, -10, -27, -32, 5, -45, -20, -1, -16, 11, -22, 18, 9, 2, -2, 33, -20, 0, -22, -35, -10, -51, -15, 4, 9, 34, -23, 16, -32, -34, 3, 17, -36, -14, -36, -8, -15, -8),
    (25, 53, -9, -13, -8, -45, 12, -4, 13, -24, -24, -13, -50, 12, -46, 10, 12, 23, 20, 37, -27, 18, -15, 8, 3, 1, -27, -19, -4, -14, -17, -4, 14, 4, 36, 37, -22, 44, -17, 5, 10, 1, -5, 0, -3, -12, 6, -13, 10, -16, 23, -24, 37, -55, -2, -5, 0, -6, -30, 25, -59, -4, -31, 38, 33, -34, 46, 27, 48, -26, 15, 8, 1, 5, -5, -18, -32, -4, -31, 21, -5, -7, 38, 33, 20, -2, 17, -26, -1, 22, -4, -16, -25, -10, -17, -1, -5, 12, -29, 6, 0, 17, -25, 8, -52, 3, 4, 30, -9, 4, -11, 21, -11, 18, -20, -16, 28, 15, 15, 3, -7, 12, 10, 24, -5, 17, -20, 18, -1, -10, 3, -18, 32, -1, 17, -1, -10, 22, -1, 25, -8, 0, -11, 12, -7),
    (10, 9, 2, -18, 1, -3, -2, -6, -15, 9, -8, 8, 20, 3, 7, 6, 20, 9, 29, -9, 38, -18, 24, -1, -4, 9, 11, -5, 13, -4, -19, 13, 20, 10, 11, 4, 11, -4, -24, -1, 3, 18, 14, 10, -14, -19, 9, 10, -4, -7, -3, 27, 35, 30, 4, 17, -33, 16, -2, 5, 12, 21, 14, 17, 27, -4, 12, 39, 56, 28, 6, 23, 7, 19, 9, -29, 18, -13, 7, 27, -4, 19, 3, 22, 5, -4, -16, 4, 23, 22, 4, -6, 7, 10, 17, 17, 11, -3, 5, 17, 36, 4, 10, 20, -23, -3, 10, -24, 29, 24, 5, 1, 28, -7, 41, 32, 53, 20, 17, 30, -6, 6, 5, -32, 16, 4, -4, 4, 5, 14, 11, 11, 19, -7, -11, -10, 24, 12, -1, -11, -4, -7, 11, 1, -5),
    (-18, 21, -16, 10, -13, 3, -29, -19, -2, 0, 19, -8, -12, -19, -16, -10, -39, 33, -28, -32, 1, -3, 8, 5, -18, 0, 8, -22, 8, -25, 0, -8, -29, 23, -17, -4, 4, -13, 8, 14, 9, 12, -10, -2, 14, -4, -5, -2, -36, 0, 25, -12, -10, -20, 13, -36, 22, 1, -5, -19, -13, -6, -33, -38, -61, 21, -41, 2, -13, 13, 6, -9, 2, 22, 14, -31, 9, -10, -5, -52, -21, 18, -29, 17, -12, 20, -14, 14, -5, 36, -13, -9, 6, -4, 21, -35, -17, -10, 16, 22, 22, 19, 25, 6, -12, 19, -55, -19, 3, -16, 19, -32, -28, 22, -20, 32, -20, 24, -25, -6, -29, 66, -20, -6, 26, 27, 28, -55, 4, -2, 4, 6, -22, 13, -33, -20, -10, 38, -11, -5, 12, 29, 12, -13, 6),
    (11, -11, 28, -37, -5, -9, -1, -16, -10, -33, -9, -16, 2, -20, -22, 17, -19, -28, -3, -35, 10, -5, -10, 4, -20, -38, -13, -23, 12, -33, -6, 15, -4, -18, -9, -2, 7, -2, -3, 15, -54, -21, -4, 6, -7, -45, 20, 2, 7, 4, -57, -32, -20, -6, 5, 22, 7, -24, -7, 0, -18, -14, 26, -2, -11, 11, -81, -14, -35, -4, -17, 32, -32, -12, -44, 36, -18, 13, 44, -17, -13, 4, -40, 19, -21, -17, -26, 11, -43, 29, -28, 16, -10, -4, 28, -5, -20, 5, -24, 1, -8, 11, -2, 28, -20, 9, 0, 11, 9, 30, 22, 13, -10, 18, -25, -17, -29, -15, -25, 12, 30, -10, -6, 48, -18, -4, 18, 5, -2, 12, -12, 4, -23, -18, -5, 12, 33, 10, -23, 17, -8, -10, 20, 5, -2),
    (36, -2, -5, 21, 37, -17, 6, -19, 20, -13, -19, -6, -28, 9, -19, 27, 6, 1, 6, 32, 20, -15, 14, -26, 4, -63, 0, -7, -45, 19, -13, -4, 11, -34, 18, 23, 0, -14, -24, 5, -18, -5, -2, -3, -29, 31, -18, -28, -8, -5, -49, -30, 19, -37, 13, -17, -9, -3, 46, 41, -23, -4, 4, 2, 18, -17, -26, 0, 18, -54, 7, 2, 13, -20, 18, 32, 13, 5, -12, 33, 30, -45, 24, -1, 15, -31, 19, 16, -37, 25, -12, 6, -22, 25, -40, -2, -4, -3, -13, -4, 27, 1, 20, 20, -24, -19, 10, 16, 18, -17, -11, 3, 3, 11, 8, -42, 17, -41, -4, -12, -14, -21, 17, -2, -11, -20, -33, 28, -20, -1, 12, -4, -12, -25, 10, -4, -5, -20, 17, -17, 1, -18, -3, 7, 7),
    (-18, -20, -15, 19, 25, 10, -3, 2, -9, 16, 4, -2, 19, -21, -15, -24, -25, -20, 30, -22, -10, 0, -16, 5, -6, 10, 27, 7, 21, -47, 20, -24, -31, -9, -5, -27, -3, -18, -22, -27, -12, 8, 20, -18, -5, -12, 18, -17, -19, -20, -23, -1, 6, 12, 4, 21, -21, -5, 28, 4, 19, -36, 33, -10, -44, -18, -30, -31, -35, -12, -21, 18, -39, 35, 25, -39, 36, -19, 17, -32, -21, -2, 10, -2, -19, -20, -7, -2, 3, 11, 1, -21, 13, -53, 15, -24, 1, 4, -20, -27, 19, -16, 6, 8, -12, -21, 2, -7, 28, 2, 27, 16, 29, 4, 10, -23, -15, -28, 1, 19, -24, 1, 14, -4, 12, 6, 36, 2, 22, -10, 23, -2, -6, -11, 9, 45, -46, 10, 12, 35, 2, -10, 20, -1, -8),
    (-9, 4, -47, -17, -5, -10, -33, 18, 5, -18, -19, 12, 7, -14, 33, 5, -12, 2, -56, 4, -38, -7, -50, 20, 0, -17, -27, 5, 11, -25, 44, 5, -4, -37, -10, 5, -18, 3, -44, 1, -36, -9, -14, -12, 4, 8, 20, 4, -19, 25, -49, -15, -43, -14, -51, 0, 52, -8, -11, 44, -5, 2, 40, 11, -13, 23, -30, -29, -50, -46, -58, 11, 53, -12, -45, 31, -12, -4, 45, 14, 7, 20, 21, 10, -26, -18, -27, 9, -1, -23, -21, 10, -11, 5, 25, 12, 4, 0, -36, -37, -34, -11, -35, 4, -8, 0, 12, 15, -8, -2, -7, 15, -9, 28, -27, -33, -12, -34, -22, 28, 26, -20, -7, 16, -29, 3, 14, 15, 9, 20, 5, -13, 2, -12, 1, -11, 21, -11, -12, 27, -6, 0, -6, 5, -6),
    (-22, 9, 2, -8, 17, -34, 18, 6, 13, 7, 19, 28, -27, 7, -8, -13, -47, -23, 19, -28, 26, -45, 7, 3, 15, 0, 24, -13, -19, -26, -19, -16, -15, -27, -2, -21, 18, -25, 6, -30, -17, -33, -7, -19, -27, -11, -2, 4, -23, 18, -19, -29, 9, -20, 7, 3, 14, -41, 44, 13, 8, 17, -39, -6, -34, 31, -39, -59, 34, -20, 28, 21, 9, -73, 54, 37, 4, -14, -13, -6, -56, -8, -46, -31, 12, -17, 12, -15, -7, -43, 34, -10, -8, -1, 6, -13, -4, 1, -1, -3, -19, -4, -6, -16, -4, -34, 34, -14, 20, 5, 12, -11, -22, 20, -13, -17, 2, -9, 4, 22, 17, -50, 58, 11, 27, 4, 8, -10, -2, 23, -57, -19, 18, -14, 1, 5, -12, -25, 16, 5, 1, -8, -7, -6, 2)
  );
  ----------------
  CONSTANT Layer_5_Columns    : NATURAL := 8;
  CONSTANT Layer_5_Rows       : NATURAL := 8;
  CONSTANT Layer_5_Strides    : NATURAL := 2;
  CONSTANT Layer_5_Activation : Activation_T := relu;
  CONSTANT Layer_5_Padding    : Padding_T := same;
  CONSTANT Layer_5_Values     : NATURAL := 24;
  CONSTANT Layer_5_Filter_X   : NATURAL := 3;
  CONSTANT Layer_5_Filter_Y   : NATURAL := 3;
  CONSTANT Layer_5_Filters    : NATURAL := 32;
  CONSTANT Layer_5_Inputs     : NATURAL := 217;
  CONSTANT Layer_5_Out_Offset : INTEGER := 6;
  CONSTANT Layer_5_Offset     : INTEGER := 0;
  CONSTANT Layer_5 : CNN_Weights_T(0 to Layer_5_Filters-1, 0 to Layer_5_Inputs-1) :=
  (
    (-29, -8, 23, 7, -15, -15, -9, 9, -7, -22, 8, -13, -5, 23, 4, -49, -11, 11, 0, 21, 14, -6, 20, -13, -35, -2, 21, -6, -11, 0, -15, -9, 2, -29, 4, -20, -33, -4, -29, -45, -34, -10, 25, 31, -14, 15, 26, -21, -29, 3, 21, -26, -10, 1, -6, -8, 8, -12, -20, 10, -38, -46, -25, -23, -22, -9, 28, 10, -28, 31, 0, -5, -7, 14, -5, 15, 19, -12, 0, -24, 30, -7, -7, 5, 28, 13, 12, 0, -46, -12, 17, 2, -7, -6, 46, 11, -27, 13, 4, 20, -2, -20, -20, -43, 27, -6, 7, -12, 18, 8, -8, -4, -26, 7, 13, 24, -20, 19, 57, 17, -50, 12, -6, -5, -23, 0, 6, -20, 14, -13, 5, 12, -17, 5, -3, -5, 12, 11, 5, 20, -9, 15, 6, 14, 2, 13, 1, -17, -3, -1, -9, 11, 7, -16, 13, -25, -5, -7, 11, -11, -19, -2, -28, -12, 11, -3, 2, 3, 0, -4, 19, -1, -13, -12, 6, -23, 1, -2, 0, 6, 4, 0, -6, -1, 2, 7, -11, 0, -5, -3, 23, 23, 11, 22, 4, -7, 0, -2, 6, -28, 6, -10, 14, 9, -7, -23, -16, -20, 2, 11, 1, -1, -7, 15, 9, 9, -6),
    (-4, 22, -38, 3, 10, -16, 7, 11, -6, -12, 12, -10, -13, -12, -4, -12, 12, -12, -11, 11, 14, 4, 6, 7, -14, 17, -43, 12, -13, -4, 7, 6, -19, -20, 34, -2, -27, 29, -4, -4, 9, 20, -20, 6, 6, 9, 18, -11, -1, -8, -32, -5, -11, 2, 17, -1, -24, -8, 44, -3, -31, 23, 22, -12, 14, -4, -20, 13, 2, 5, 20, -6, -1, -7, -17, -20, -37, -18, 15, 7, -18, 4, 12, 31, -23, 11, 19, -5, -6, 2, -14, -35, 27, -1, -27, 19, 10, -7, -6, -11, -38, -28, 29, -12, -6, 21, 20, 39, -22, 33, 47, -35, -6, -4, -3, -55, 20, -10, -53, -3, -8, 5, 8, -15, 4, -26, 12, -27, 16, 36, -16, 29, -12, 22, 34, -16, 10, -8, 25, -46, 0, -9, -20, -15, -1, -5, 5, -18, -2, 7, 18, -5, 2, 24, 1, 4, 35, 3, 12, 21, 19, -16, 12, -20, 10, -20, -12, -19, -1, -7, 0, -8, -7, 39, 3, 4, 1, 22, -5, 6, 23, 3, 21, 32, 2, -21, 13, -22, 10, 5, -8, -31, 3, -22, 22, -12, -20, 24, -9, 21, -18, 8, -5, -14, 22, -15, -2, 19, 10, 12, -2, -21, 0, 3, -4, -18, -3),
    (8, -12, 50, -12, -6, -32, 13, -50, 26, 30, -12, -2, -40, -2, 33, 11, -30, -12, 37, -5, -13, -8, -5, 3, 21, -15, 20, -17, 6, -48, 3, -7, 21, 34, -37, 25, -9, -5, 12, 23, -27, 10, 23, -5, -5, -1, -11, 7, 35, -18, -17, -20, 16, -27, -4, 13, 27, 21, -27, 18, 11, -36, -5, -16, -8, -4, 2, -15, -1, -12, -13, 3, 32, -19, 25, -15, -2, 6, 0, -36, 28, -14, -47, -35, -8, -30, -18, -31, -36, 13, 14, 14, -26, 18, 4, -42, 38, -15, 33, -23, 15, -22, -12, 6, 19, -22, -50, -30, 15, -39, -32, 21, -19, -10, 27, 12, -3, 11, 6, -19, 19, 9, -5, -28, 36, -32, -8, 25, 1, -23, -24, -19, -12, -22, -24, -9, 2, 4, 0, -7, 12, 13, -3, 6, -30, -4, -11, 21, 9, 20, -9, -5, 0, -22, 11, -33, -5, 28, -20, 20, -3, 37, 4, 12, -17, 11, 10, -29, 14, 12, 2, 5, 6, 34, -14, -4, -11, -18, 11, -28, 19, 44, -20, 19, 10, -5, -1, 22, 6, 24, 16, -25, 3, 12, -25, -1, 4, 22, 0, -19, -5, -9, -10, -8, 1, 26, -3, 18, 1, -1, 4, 20, 4, 10, 15, -13, -1),
    (-13, 24, -22, -4, -6, 5, 2, 1, -8, -26, 1, -18, -6, 22, -14, -6, -9, 16, -13, 11, 4, 19, 12, 1, 9, 7, -3, -22, -19, 12, 7, 6, -22, -44, 1, -17, -5, -6, -15, -8, -13, 2, -15, 17, -9, 30, 16, -14, 30, -3, 13, -22, -3, -7, -4, 14, -4, -2, -10, 4, 1, -29, 0, -22, -7, -6, -10, -2, 2, 20, -20, 6, 5, 18, -23, 24, 19, 1, -12, -16, -11, -17, 5, -12, -6, 21, -29, -1, -2, 27, -12, 30, -13, 12, 18, -4, -1, 7, -28, 35, 13, 25, -14, -11, -20, -37, 1, -29, -19, 52, -44, -6, -15, 15, -16, 43, -33, 22, 36, -41, 20, 17, -31, -2, 0, 20, -11, 4, -13, -15, 9, -8, 2, 20, -21, -29, -4, 3, -26, 14, -28, 20, 11, -37, 6, -8, -2, 19, 12, -24, -1, -13, 20, 11, -6, -5, -29, 2, 2, -19, -16, -25, 27, -20, -24, -28, -14, 24, 4, 16, -2, 22, 37, -38, -23, -16, 19, 10, -7, -12, -22, 0, -3, -21, -34, -10, 18, -3, -25, -43, -2, 10, 2, -7, 16, 13, 28, -19, -33, 4, 9, 26, -12, -2, -28, 18, 1, -5, -28, -19, -32, 1, -7, -35, 4, -1, -5),
    (-16, 6, 21, -10, -19, 0, -18, -18, -27, -25, -5, 35, 52, 16, 20, 34, 26, -32, 12, 7, 37, -19, 12, -19, -4, -10, 26, -25, 3, -15, -6, -20, -7, -8, 16, -13, 33, -12, 17, -7, -27, -22, 16, 11, 20, -1, 1, -6, 13, -6, 6, -18, -9, -58, 4, -8, 1, -18, 4, -4, 1, -27, 11, -13, -53, -19, 14, -3, -16, 1, 20, 11, 0, -18, 37, 1, -2, -33, 4, -3, -13, 24, 13, -4, 24, -28, 39, -23, -2, -21, 25, 12, 4, -23, 6, -24, 27, -34, 29, -7, 22, -29, 0, 16, -2, 29, -10, 2, -22, -26, -5, -30, -45, -17, 43, 9, -14, -4, 5, -7, 11, -24, 12, 3, 24, -8, -14, 25, 20, 8, 4, 2, -3, -47, -22, -13, -44, 7, 16, 12, -26, 6, 19, -6, 21, -35, 26, -2, 23, -9, 30, -2, 5, 18, -13, -5, -16, -34, -19, -5, -20, -1, 18, 5, -33, 4, -11, 9, -3, -18, 31, -8, 20, 18, -6, 9, 26, 15, -20, -20, -12, 7, -26, -6, -20, 11, 28, 23, -21, 16, 2, -5, -6, -4, 14, 1, 16, 13, -15, 22, 15, 6, 6, -9, 19, 12, -39, 19, 6, 14, 16, 21, 13, -10, 5, -10, 15),
    (-10, -26, 2, -44, -29, -12, -80, -14, -29, 34, -1, -26, 3, 20, 18, -2, 20, -45, -4, -24, 17, -4, -14, -52, -18, -12, -12, -27, -31, -23, -39, -5, -35, 30, -34, -69, 23, 13, 7, 28, 10, -21, -12, 20, 15, -5, -5, -33, -23, -9, 16, -23, -29, -22, -27, -1, -29, 3, -28, -62, 21, 36, 1, 36, 3, 0, -8, 17, 24, 10, -5, -42, -4, 28, -30, 5, 11, -7, -20, 7, 13, -15, 6, 13, 39, 22, -13, -1, 21, 18, -16, 12, -4, 4, -13, 1, -33, 20, -43, 6, 11, 0, -6, -25, -4, 26, 5, 25, 36, 50, 3, 5, 36, 24, -29, 20, 13, 4, -10, 32, -29, 9, -12, -2, -3, 21, 11, -26, -30, 0, 5, 1, -6, 3, 21, -20, 16, 9, -20, 36, 12, 13, 6, 24, 3, 5, -23, -28, 10, -3, -2, -11, -13, 13, 6, -16, -1, 0, 5, -3, -20, -10, -13, 7, 4, 12, 11, -1, -9, -2, -34, -29, 19, 3, 3, -32, 12, 29, -12, -7, 3, 4, 15, -4, -31, -11, -12, -5, -19, 14, 18, 16, 30, -5, -16, 0, 21, -6, 4, -19, 24, 28, -20, -11, -1, -7, 18, -21, -38, -3, 5, -22, -38, 9, 10, 7, -2),
    (11, -43, 29, -23, -18, -14, -38, -7, -22, -33, -14, 2, -2, 0, 9, -4, -28, -35, -16, -11, -5, -13, -6, -42, -7, -21, 3, 9, -17, 6, -27, -2, -40, -40, 3, 4, -10, 16, 35, 8, -23, -28, -19, -11, -8, -26, -6, -31, -14, -12, 24, 11, -5, -3, 5, 25, -72, -29, 23, -4, -20, 6, 12, -15, -1, 4, -14, 5, 20, 10, -2, -9, -26, 20, -35, 40, -23, -9, -19, 14, 11, -12, 0, 2, 36, 32, 45, 3, 28, 3, 4, 5, 7, -13, -12, -1, -18, -10, -38, 24, -16, -26, -29, 10, -1, -20, 1, -22, 27, 22, 26, 26, 21, -10, -15, 2, 3, 9, -5, 6, -12, -28, 0, 5, -25, -6, -12, 24, -34, 9, 23, 4, 12, 15, 45, -4, -6, -11, -31, -5, 11, -20, -18, -16, -22, 26, -36, -20, 4, -16, 12, -6, 9, 15, 7, 22, 12, -22, 28, -5, 5, -7, -5, -6, 0, -5, -19, 32, -42, 32, -37, 1, 12, -38, 9, 7, -10, 34, 0, 27, 24, 0, 31, -18, 11, -3, -14, -4, 27, 2, -14, 42, -39, 11, -10, 17, -24, -32, 16, 2, -29, 8, 15, 7, 21, 25, 34, -18, 11, -9, -25, 14, 17, 10, 0, 18, 1),
    (17, 1, -23, -27, -12, 10, 27, 8, 15, 10, 21, 24, 9, -4, 1, 33, 4, 4, 23, -7, 13, 10, -11, -21, 3, 4, 19, -49, -16, 3, 15, -23, -23, 20, 10, -3, 24, -13, 14, 23, 12, -24, -24, -8, -16, 15, -8, 12, -7, -2, 32, -2, -24, 5, 26, -17, -32, -31, 14, 7, -8, -15, -10, 3, 8, 8, -1, 2, 0, 21, -5, 3, 46, -12, -8, -26, -11, 20, -14, 28, -13, 4, 1, 5, 16, 25, -17, 22, 7, -2, -15, -5, -2, -4, -17, 3, 18, -20, -12, -35, -21, 3, 15, -5, -70, -23, 32, 13, 8, 21, 42, 14, 20, -26, -47, -19, 35, 6, -44, 30, 8, 17, -20, 2, -21, -3, 29, -17, -30, -26, 15, 24, -14, -4, -12, 0, 23, 21, -20, -8, 15, -4, -16, 5, 23, -5, -31, -18, 11, 14, 3, 6, -19, -24, 25, 3, -2, 39, 19, 6, 6, -22, -26, -5, -14, -6, -33, -5, 20, 1, -31, -16, -3, -20, 9, 6, -45, -9, 23, 21, 5, 10, 9, 8, 7, 6, -34, -19, 8, -12, -26, 11, 15, 20, -24, -9, 6, -8, 3, -7, -14, -16, 6, 23, -7, -11, 1, -1, 23, 22, -20, -4, 11, 1, -12, 0, -2),
    (2, -24, 51, -6, -14, -33, -5, -40, -13, -37, 13, -19, -25, 43, 1, -21, -2, -34, 10, -11, -1, 5, -22, -20, 11, -9, 41, 8, -6, 1, -1, -38, -3, 22, 5, -22, -16, -39, 3, -28, -13, 2, 36, -6, -27, -3, -26, -14, -24, -9, -8, -8, -32, 17, -6, 11, 12, 2, -11, -5, 19, -23, 27, 26, 13, -27, 0, 3, -5, -22, -25, -15, 23, -20, 38, 12, -26, 36, 9, -24, 20, 15, -5, -9, -38, 6, -19, -5, -4, 19, 4, 21, -15, 27, 2, -24, 45, -49, 66, 6, -20, 28, 19, -42, 34, 21, -9, -27, -36, -32, 12, 14, -13, -11, 32, 16, -54, 18, -19, -35, 28, -20, 0, -1, 2, 11, 14, -2, 31, 39, -24, 4, 2, -32, 15, 12, -6, 3, 37, -4, -26, 4, -33, -30, -12, 0, 27, 12, -31, 2, -4, 3, 17, 0, -1, 4, -1, 16, -21, 3, -20, 5, 11, 7, 9, 5, 2, -8, 14, -11, 46, 12, -17, 4, -11, 9, 18, -13, -6, -6, -20, 37, -19, 3, -20, 5, 2, 9, -10, 13, 8, -21, -13, -4, 14, -8, 4, 4, 4, 12, 4, -18, -11, -12, 19, 5, 17, -10, -18, -12, -1, -12, -3, 19, 5, -2, 0),
    (-17, 11, 3, -23, 22, 3, 6, -3, -2, -13, -5, -13, -1, -27, 3, 7, -16, -9, -20, -11, -22, 30, 20, -1, -37, 6, 3, -29, 20, -1, 11, -3, -1, -27, 6, -20, -5, -48, -25, 23, -28, 3, -29, -1, -2, 20, 22, 12, -33, 2, 4, -24, 14, -9, 15, -12, -4, -15, -7, -9, -26, 4, -14, -17, -22, 12, -18, 10, -7, 8, 4, 10, -7, -1, 6, -11, -27, 32, -13, 0, -39, -12, 27, -21, 7, 42, -18, 27, 1, -19, -26, 4, 11, 34, 20, -22, -36, -3, 3, -10, -39, 35, 21, -27, -39, -5, 52, -12, 24, 45, 23, 35, 9, -14, -38, 10, 7, 40, 21, -12, -13, 13, -7, -12, -17, 12, 28, -31, -19, 8, 36, -10, 17, 21, 37, 0, -7, -9, -8, 18, -3, 4, 14, -4, 9, 12, -3, 1, -10, -19, -5, -9, 14, 5, 0, 36, 0, 15, -35, -4, 9, 1, 6, -22, 9, -15, -29, -4, 1, 2, 2, -12, -13, -7, -4, -21, 10, 27, -12, 48, 2, -1, 21, -3, 2, -14, 10, -24, 28, -16, -24, -6, 12, -14, 4, -6, -10, -13, 2, -7, 20, 29, -17, -1, 12, -13, 20, 4, -4, -28, 12, -13, 15, -10, -22, -6, -8),
    (-30, -8, -1, -21, -22, -21, 9, -8, -52, 5, 10, -7, 3, -29, 6, -19, -9, 13, -28, -19, 4, -4, -2, 34, -43, 6, -5, -3, -31, -29, -16, -10, -70, -28, 43, 15, -12, 21, 35, -21, -16, -4, -8, -37, -6, 0, -14, -15, -2, 27, -8, -6, 4, -31, 4, 7, -5, 1, -4, -6, -35, 9, 20, -25, -18, -10, -37, -44, -9, -38, 2, -47, -2, 23, -30, -8, -25, 5, 12, 4, -50, 13, 5, -3, 39, -6, 19, 3, 49, -28, -41, -8, 12, 10, -2, 4, -37, 10, -12, -13, -31, -2, -9, -20, -12, 29, -29, -29, 29, 25, 30, 39, 33, -24, -5, 0, -6, -8, -2, -10, -62, -26, 6, -15, -37, -12, -17, 4, -10, 27, -54, -35, 16, 6, 26, 21, 12, -29, 6, -4, -3, 17, 4, -19, -17, 27, 4, 3, -2, 5, -10, -20, 30, 29, -9, 15, -4, 12, 24, 5, -29, -22, 17, 9, -32, -8, 9, 14, -8, 11, 1, 23, 7, 5, 0, -6, 16, -12, -20, 3, 41, 21, 8, 4, 5, -17, 19, 28, 0, -2, 0, 4, -5, 19, -6, 12, 26, 29, 5, -3, -12, -13, -12, -8, 45, 43, -2, -8, 3, 9, 24, 21, 15, 3, 3, 4, -1),
    (-20, 7, -70, 1, 4, 2, 0, 21, 0, -20, 19, 11, 0, 15, 0, 5, 33, 11, 3, 13, 20, -6, -6, 12, -17, 2, -25, -16, -57, -23, 17, -2, -40, -20, 22, 20, -4, -3, 10, -8, 40, 4, -54, -13, 36, -11, 5, 42, 5, -28, 36, -17, -6, -11, -20, -32, -14, 28, -4, -14, -16, -12, -5, 8, -11, 9, 5, 4, 2, -2, -25, 13, -18, 10, -18, -7, 12, 0, 19, 3, 14, 0, -11, 13, 7, -25, -3, 8, 11, 3, -7, 4, 20, 2, 0, 35, -43, 15, -33, -18, -26, -26, 23, -16, -48, 10, 24, 29, 29, -14, 12, -11, 6, -13, -67, -12, 9, 5, -10, 40, -27, -16, 13, -18, -1, -24, 23, -27, -19, 34, -37, -11, -10, -5, 49, 1, -58, -6, -19, -35, -27, -5, -19, 19, 0, -5, -11, -10, 11, 5, -1, -4, 5, -3, 20, 18, 6, 6, -2, -2, 2, -27, -6, 4, -18, 12, 5, 3, -22, 12, -13, -9, -9, 9, 8, -8, -6, 29, 12, 16, 40, 8, 10, 19, 24, -16, -23, 18, -13, 1, 7, -13, -3, 20, -12, -7, -4, 1, -26, -9, -16, -13, -14, 11, 16, 12, 2, 17, 16, 4, -45, 7, -7, 18, -13, -12, 12),
    (2, -15, -21, -16, 1, 5, -1, -6, -2, 20, 16, 19, 14, -13, 28, 12, 3, -6, -27, -25, -9, -11, 7, 4, -15, -18, 11, -12, 22, -15, 1, -37, -21, 5, 21, 9, 3, -15, 20, -15, -6, -3, -30, -13, 27, -3, 9, 26, 21, -23, 0, -8, 6, -4, -9, -7, 4, 19, 17, 1, 0, -9, -13, -23, 11, 18, -13, 9, -3, -13, -10, 24, 0, -8, 5, -25, 9, -19, -14, -41, -51, -6, 12, -2, 15, 14, 28, -16, -28, -29, -20, -37, 7, -25, 1, -10, -6, -20, 6, 43, 26, -28, 13, -6, -12, 54, 19, -4, -18, 10, 12, -68, -4, -8, -1, -11, 10, -21, 13, 12, 4, -7, 20, 12, 36, -1, 4, 4, 3, 40, 14, -15, -1, 4, 19, -29, 4, -12, 3, 1, -4, -20, -6, 9, -23, -13, -19, -18, -2, -6, -50, 19, 9, -10, 9, -7, 7, 21, -37, -17, 19, -28, 3, 14, -10, -12, -16, 3, -5, -7, -2, 28, 5, -23, 21, 22, 4, 38, 7, 4, 34, -19, 34, -3, -2, -16, 15, -3, -25, -50, 1, 6, -5, -28, 13, 35, 26, 4, 22, 6, 6, 34, -8, -8, 18, 0, 28, -11, -27, 2, -6, 3, -12, -45, 13, 4, 29),
    (24, 19, 0, -28, -21, 26, -1, 10, -3, -27, -12, -4, 22, 23, -4, 17, 26, 2, -45, -13, -16, 14, -3, 2, 19, 8, -5, -27, -20, -9, 28, -25, -29, -50, 31, 1, -11, 14, -46, -9, 9, -1, -24, -1, 10, 8, -17, 14, -2, 16, 6, 12, 14, -12, 28, -14, -12, 1, 29, 3, -13, -3, 5, -15, -7, 25, -14, -5, -12, -9, -1, 12, 12, -2, -28, -53, -20, 17, -9, -9, -30, -5, 16, 6, 24, 11, 14, 28, 31, -21, -50, -24, 30, 11, -23, -16, 11, 8, -34, -12, -40, -12, 34, -13, -46, -27, 37, 40, -11, -22, 7, -13, 28, 21, -65, 5, 18, 3, -9, 7, -6, 5, -11, -1, -5, -9, 35, 4, -21, -9, 25, 5, -12, -1, 39, -21, -1, 14, -17, 14, -15, -4, 19, 10, 29, -13, -8, -27, -3, -1, -9, -9, -28, 22, 9, 18, 20, -4, 4, 12, 5, -35, -26, 3, 17, -4, -23, -18, -9, 17, -34, -12, -14, 4, 20, 3, -19, 1, 6, 18, -4, -28, 12, 3, 30, 18, -22, 13, 16, 10, -5, -5, -10, 11, 9, -2, -7, -9, 20, -7, -2, 9, 6, -5, -13, -11, 9, 2, -2, 18, 21, 12, -4, -9, 8, -8, -1),
    (14, -27, 25, -14, 13, 19, -9, -2, 20, 13, -16, -28, -19, -18, -20, 2, -27, 19, 36, 10, -34, 12, -13, -31, 46, -21, 12, 14, 20, 35, -18, 38, 31, -4, -10, -28, -5, -12, -60, 18, -4, 29, 55, 3, -15, -15, -7, -48, 44, 2, -19, 11, 12, 39, -16, 25, 12, -22, -7, -7, 13, -7, -30, 32, 17, -8, 10, 8, 2, 20, -12, -24, -8, -11, -11, 45, 12, 8, 4, 17, 9, -6, 7, -12, -23, -9, -1, -27, -5, 28, -1, 7, -6, -4, -10, -10, 3, -20, -37, 44, 7, -5, -13, 23, -5, -27, 27, -20, -13, 7, -22, -7, 7, 12, -24, -3, 24, -18, -16, -8, 3, -7, -23, 11, -3, -14, 11, 12, -52, -39, 34, 5, -18, 8, 17, -8, 19, 6, -44, -24, 18, -26, -9, 11, 18, -6, -7, 4, -13, 2, 0, -1, -29, -1, 20, -7, -21, -12, 6, 6, 4, -11, -18, -11, 13, -18, -19, 22, 1, 1, -15, -11, -11, 6, 28, -15, -34, 2, 19, 21, -16, 14, 30, 21, 20, 12, -27, -18, 2, -8, -20, 20, -4, -20, 13, -29, -23, 20, 28, -38, -14, 19, -13, 29, 18, 9, 29, 20, 5, -20, 15, 0, -1, 10, 2, 5, -3),
    (7, 30, -44, -4, -9, 6, 5, 10, -4, -13, -2, 17, 17, -8, 28, 33, 29, 4, -29, -10, 17, 5, -23, 12, -11, 13, -16, 13, -15, -3, 25, 10, -28, -12, 6, 13, -3, 35, 11, 11, 19, 24, -40, -9, -5, 10, -6, 13, 4, -3, -19, 8, 16, 2, 11, -11, -15, -12, 27, 2, -14, 19, 5, -9, -7, 5, -5, -8, -1, 4, 7, 31, -4, 18, -53, 3, -10, 11, 20, 11, 3, -25, 17, 23, -19, -2, 0, 11, 39, 7, -20, 0, 12, 21, -30, 25, -9, 36, -20, 20, -11, -11, 9, 1, 5, -21, -14, 10, -19, 19, 1, 1, 33, 7, -8, -7, 5, -7, -18, 53, 16, 20, 5, 20, -4, 13, -4, -8, 5, -11, -7, -26, -11, 12, -14, 3, 2, 30, 1, 5, -12, 3, 3, 6, -13, 17, -23, 5, 0, 22, 8, -17, -10, -9, 0, -3, 4, -13, -10, -1, 6, 15, 1, 12, -2, 23, -6, -2, -2, 28, -20, -3, -5, 12, -18, 0, 9, -22, -12, 29, 2, -13, -16, -10, 12, -1, -6, 11, -12, 12, -4, -6, 16, 23, 8, -7, -2, 13, 0, -16, -3, 0, 1, 0, 16, 12, -9, 28, 5, 28, 12, 21, -17, 8, 13, -7, 3),
    (2, 20, -36, -12, 5, -11, -1, -11, 21, 6, 10, 21, 11, 0, 0, -18, 44, 15, -19, 2, -1, 0, -13, 12, 3, 11, -45, 10, 3, 5, 9, -10, 20, 18, 0, 28, -5, 12, 20, -38, 26, 11, -10, 0, -18, -2, -1, 30, 24, -17, -5, 27, 8, 9, 14, 7, 4, 0, -19, -17, -2, 0, 11, -8, 1, -9, -29, -8, -11, -4, 4, 19, -7, 2, -58, -20, 24, 12, 17, -35, 23, 46, 5, -4, 1, 5, 24, -19, -14, 8, -1, -19, -29, 4, 9, -17, 0, -16, -43, 16, 18, 4, 13, -35, 30, 43, -13, 1, -2, -4, 26, -29, -11, -20, -23, -21, -34, 5, 11, 7, 25, -12, -22, 28, 32, -12, 10, -12, 6, 22, -42, -61, -14, -6, 4, -23, -40, -3, 5, -31, -42, 8, 21, -10, -10, -11, 17, -19, 13, 5, 4, -11, -10, 12, -3, -10, -7, -6, 23, 5, -6, -7, 11, -9, -28, 3, 12, -41, 3, -21, 21, -11, 43, 15, 4, 17, 5, 5, -18, -25, -21, -8, 0, -15, -13, -15, 16, -41, -49, -2, 11, -14, -2, -38, 2, 6, 30, 4, 18, 29, -20, 17, -6, -22, -20, 14, -7, -33, 1, -3, -14, -37, -20, -24, -2, 12, -5),
    (4, -16, -9, 5, 29, -5, -5, 0, 30, 26, -12, 7, -7, -6, -3, -4, 6, -35, 6, -15, 17, -19, -11, 22, 27, -40, -6, 13, 19, 8, 5, 13, 28, 56, -15, 15, 5, -31, 13, 2, 11, -21, 4, -31, 17, 18, -38, 42, 23, -2, -4, -1, -2, -3, -13, 9, 17, 50, 6, 10, -3, 6, 7, 11, -1, 1, 6, -17, 28, -3, -35, 29, -9, -4, 20, -8, -32, -7, -24, -25, -10, -16, 14, 10, 16, 20, -43, 10, 12, -11, 3, -11, 7, 5, -35, -5, 15, 7, 3, 7, -20, -8, -8, 15, 20, -30, 3, 35, 10, 13, -25, 20, 19, 2, 4, -3, 4, -4, -55, -27, 12, 16, -16, -16, 20, -22, -4, 10, 12, 11, -4, 46, 24, 17, -1, -7, 20, 1, 18, -6, 20, -19, -39, 1, 24, -19, 29, -15, -28, 3, 7, -24, 29, 25, -7, 8, -3, 10, -5, 1, 6, 8, 28, 20, -10, 25, -9, -19, 25, -36, 47, -12, -5, 5, 29, -24, 28, 20, -9, 11, 14, -21, 15, 20, -12, -12, 50, -8, -20, -5, -13, -35, 23, -21, -18, -13, 4, 6, 12, -8, 29, 23, -3, 17, 24, -1, 20, 19, -14, -5, 19, -15, -3, -16, -28, -5, 4),
    (-31, 2, 1, -10, 6, 2, 26, -3, -3, 3, 10, -5, 13, 2, 25, -4, -43, -6, 22, -21, 0, 6, -9, 19, 38, -4, 11, -4, 6, -35, -18, -17, 4, 18, -6, -5, 0, 13, -8, -69, -40, -16, 8, 10, -29, -24, 8, -4, -6, 11, -4, 21, 32, -5, -35, 6, 7, -15, 4, -12, 18, -12, -31, 4, -7, -5, -5, 9, 7, 18, 13, -5, -47, -2, 33, -3, 28, -20, -10, -40, 27, 15, 9, -14, 8, 31, -4, -25, -64, -27, 25, -5, -1, -6, 10, 2, -10, -9, -12, 20, 40, -7, -33, 8, 22, 6, -4, -23, 14, 4, -33, -34, -47, -15, 4, 7, -32, 10, 39, -1, -21, -9, -22, 19, 21, 0, -8, 9, -15, -16, 12, -19, 11, 4, -11, -4, -7, -1, -12, 24, -11, 0, 27, 1, -44, -7, 22, 3, 10, -25, -14, -18, 16, -11, 2, -19, -16, 11, 1, -37, -41, -11, 35, 6, -34, -11, 4, -2, -45, 6, -3, 26, 12, -3, -19, 17, 19, -12, 12, -18, 12, 18, -18, -19, -32, -11, -2, 5, -12, 20, 36, -11, -8, -1, -13, 8, -8, -5, 3, -5, -5, 13, 20, -20, 15, 4, 15, -4, -29, -2, -11, 5, 0, -12, 20, 7, 2),
    (12, 7, 9, 21, 13, 12, 3, -7, -6, 0, -6, -14, 17, 5, -21, 24, -5, 4, 17, 20, 2, 3, 22, 29, 5, 20, 36, 16, -4, 22, -6, -5, -11, -22, 20, -36, 44, 41, -21, 28, 7, -13, -4, 28, 0, 4, 21, -8, -9, 10, 33, -5, -5, 17, -9, 1, -2, 4, 17, -11, 15, 20, 7, -5, 3, 1, 10, -1, -4, -9, 6, -16, 7, -36, 29, -11, -22, -37, -43, -37, 11, 34, -20, 1, -7, 32, -17, -24, -9, -21, -26, -13, 5, -24, -28, -25, -20, 0, 27, -21, -40, -23, -34, -12, -17, 12, -8, 1, -5, 20, 15, 7, -2, -20, 10, -2, 19, -6, -16, -7, 4, -20, 18, -26, -51, -27, -15, -2, 5, 22, -32, 1, 14, 9, 10, 27, -3, -28, 6, 15, 8, 2, -21, -4, -3, 12, -10, -18, 11, 14, -22, -20, 4, -11, -13, -13, -12, -30, -22, 7, 18, 4, 31, 37, -30, -2, 0, -9, 42, 13, 5, -32, 21, 14, -28, 29, 31, -28, -68, -4, 9, -15, -10, 21, 5, -2, 43, 11, -7, 24, 8, -13, 42, -10, 24, 4, 29, -23, -6, 12, 14, 5, -47, 3, 29, -27, -11, -13, -5, 0, 30, 21, 5, 24, 3, 6, -1),
    (22, -12, 13, -20, 7, 25, -7, 22, 17, -39, 7, 29, -3, -16, -19, 12, -13, 5, 1, -16, 4, 3, -9, -20, 17, -4, -3, -54, -46, -11, -33, 22, 4, -34, -5, 41, -11, -24, -6, -17, -17, -5, -6, -9, 9, -6, -25, -13, 9, -27, -3, -42, -29, 7, -21, -6, -14, -20, -25, -7, 7, 3, 9, -5, -3, -12, 5, -35, 28, -19, -37, 16, 18, -4, 3, -13, 33, 36, 4, 31, 12, -19, -14, -18, 24, 21, -21, 44, 1, 17, 26, -4, 2, -11, -3, -32, 36, 18, -14, -30, 37, 42, -20, 32, 44, -13, -15, 13, 26, 9, -15, 46, 28, 21, 35, -11, 17, -12, -34, -39, 12, -2, -20, -20, -14, 7, -13, -4, -5, -17, -5, -2, 5, -7, 25, 8, 16, 2, -29, -2, 14, -12, -14, -11, 34, 19, 5, 6, 35, 5, -2, 10, 13, 6, -4, 9, 22, -1, 0, 3, 12, 12, 16, -6, 3, -14, -7, -21, 15, 18, -51, 1, 21, 8, 3, 23, 12, 13, -4, 24, 32, 13, -14, 13, 29, 17, 4, -5, 19, -27, -28, -25, 18, 8, 5, -20, 14, -3, -3, 5, 7, 19, -13, 15, 18, 2, 12, -6, 15, 7, 18, -4, 12, -24, -25, 13, 0),
    (10, -28, 13, -15, -16, 1, -47, -20, -10, -12, 13, -7, 11, 43, 1, 22, -4, -34, -10, -15, 8, -28, -23, -36, -8, -11, -10, -18, 39, -5, -44, -10, 14, -10, -10, -15, 17, -20, 10, -22, -2, -10, -4, 15, -11, -12, 5, -14, -9, 19, -35, -7, -3, -11, 1, 14, 6, -16, -27, 11, 21, -31, -11, -23, 16, -7, 13, 0, -12, -9, 9, 6, -1, 9, -20, 15, 27, 17, -21, 19, 14, 3, -46, -13, 14, 3, -36, -40, -3, 10, 31, 23, -25, -12, 16, -34, -13, 14, -32, 30, 37, -7, -35, 45, 20, -14, -4, -28, 3, -20, -10, -4, 20, -3, 13, 25, -4, -29, 15, -7, 13, 19, -3, -1, 23, -5, -9, 24, 2, -19, 4, -21, 13, -23, 3, 7, 5, -4, -1, 12, 22, -8, -2, 9, -25, -10, 7, 29, 20, -20, -5, -5, 25, -13, 3, 10, -71, -12, 3, -15, -8, 21, 11, -14, -19, -7, 9, 3, -11, -3, -38, 17, 3, -3, -10, 18, -12, -19, 16, -4, -6, -21, 8, -2, 13, 2, -4, 6, -4, 5, 2, 3, 18, 4, 12, -18, -23, -21, 23, 5, -24, -13, 11, 3, -3, 10, 13, 14, 8, -4, -14, -22, 24, -14, -18, 12, -3),
    (20, -2, 4, -3, 9, -21, -5, -24, -2, -11, 2, -8, -11, -38, 1, -32, 7, 2, 4, 1, 18, -10, -7, 5, 5, 7, 0, -9, 13, -29, 5, -1, -1, -28, 1, 5, 3, -53, 7, -25, -3, 12, -3, -10, 19, -1, -8, 10, -11, 4, -40, 5, 6, -4, 12, 0, 0, -29, 12, 30, -10, -25, 4, -62, -3, 4, -13, -13, 11, 5, -7, 10, 19, -6, -6, 7, 1, 41, 6, 23, 9, 4, 13, -13, 15, -4, 1, 32, 11, 5, 40, 5, 9, -14, 3, -11, 22, -10, -16, -10, -19, 24, 10, 24, -4, 4, 38, 11, 42, -4, 33, 58, 35, -15, 51, 13, 30, -6, 4, -36, 24, 12, 1, -23, -33, 5, 9, 6, -9, 13, 25, 13, 15, 2, 29, 17, 27, -8, -18, 6, -8, -9, 4, -38, -19, 4, 10, -5, -28, -44, -12, -8, -25, -20, 5, -32, -26, 8, 1, -1, -4, 1, -22, 12, 2, 9, 14, 1, -5, -20, -10, 14, -31, -33, -36, -10, -34, -36, -2, -31, 11, 44, -8, 16, 2, -19, -18, 18, 15, -11, 6, 16, -30, -25, -1, 0, -61, -36, -25, -6, -35, -37, -32, -8, 18, -7, 8, -1, -30, -26, -3, 20, -10, 14, -3, 30, -1),
    (-13, 6, -4, 11, 12, -22, 6, 5, -13, -35, 4, 4, -25, -16, -12, 9, -9, 6, 1, 32, 2, -13, 15, -2, -22, -4, -31, 13, 20, -6, -23, 12, 4, -32, -5, -8, 7, -17, -52, 2, -20, 6, 29, 28, -33, -9, 31, -37, 3, 7, -18, 18, -5, -4, -4, 6, -12, -20, -31, 18, 26, -7, -2, -7, 7, -11, -55, -24, -12, -15, -5, -21, -10, 6, -1, 9, 14, -18, -3, 34, -18, -15, 5, -4, 17, -35, -8, 12, -2, 12, 38, 28, 13, -20, 9, -24, -4, 8, -7, 26, -5, -12, 2, 33, -45, -26, 4, 3, 0, -27, 11, 20, 8, 11, -4, 8, 10, -24, -4, -28, -26, -4, 27, -4, -44, -17, 3, -12, -19, 13, -44, 29, -1, 16, 29, -17, 6, 0, -3, -13, 15, 12, -27, 23, 5, 25, -37, -2, -16, 9, 15, -3, -10, -20, 12, 9, 14, -3, 0, 3, 23, 4, -26, 4, 11, 0, -25, -7, -24, -9, 16, -49, -23, 0, 20, -20, -5, 2, -19, 10, -3, 0, 11, 11, 17, -16, 11, -29, 23, 7, -39, 20, -11, -13, 8, -44, -6, 29, -21, -46, 33, 14, -19, 28, -1, -15, 4, 3, -9, -22, 19, 17, -17, -11, -5, -12, 9),
    (10, 1, -34, -2, -4, 12, -13, -3, 8, -5, 12, 27, 11, 22, -4, -12, -2, 4, -13, 6, -8, 7, 13, -7, -6, 12, -38, 4, 20, 4, -18, -24, 17, 11, 3, 25, -11, 36, -4, -28, 19, 8, -46, 4, -31, 20, 3, -43, -5, 10, -34, 8, 16, 11, -4, -19, 10, -2, -12, 20, -6, 25, 4, -33, 21, -2, -23, 8, -22, 20, -5, -26, 41, -13, -28, -32, 20, -31, 2, -26, 4, 49, -5, 8, 4, -21, 2, -2, 6, -5, 9, -43, -8, -26, -20, -4, 24, 16, -8, 2, 31, -31, -24, -28, 32, 77, -21, 25, -27, 5, 17, -27, 2, 8, 11, -47, -33, -13, -17, -9, -25, 13, 13, 25, 32, 5, -28, -1, 44, 27, -19, 14, -30, 16, -1, -29, -33, 8, -18, -13, -18, -22, -15, -20, 9, -19, -9, -5, 34, 5, 24, 25, 2, 17, -14, -1, 11, -38, 6, -6, 12, -16, 8, -13, -4, -25, 4, 0, -4, -18, 10, -10, 27, -15, 12, 33, 7, 31, -12, -14, 8, -36, 0, 14, -5, -14, 27, -28, 9, -38, -6, 14, 14, -19, 8, 2, 23, -8, -3, 21, 9, 18, -23, -41, -7, -29, -9, 9, -35, -17, 23, -35, 14, -39, 14, 20, -5),
    (-12, -45, 19, 20, 5, 13, 0, -10, -8, 12, 2, 0, -4, 4, 22, -17, -21, -35, -6, 4, 32, -12, -8, 27, -4, -19, 28, -25, -8, -9, 6, -9, -30, 25, -18, -1, -7, -15, 1, 8, 12, -10, 8, 4, 9, 8, -13, 36, 6, 2, -2, -7, -1, -18, 19, -18, 2, 11, -7, -15, 31, 12, 10, 10, 24, -20, 4, 10, -4, 21, -23, 13, -22, -45, 34, -2, -44, 4, -1, 0, -17, -33, -12, -29, -3, 4, 0, 17, 1, -16, -2, 6, 18, 20, -11, 21, -16, -24, 34, -4, -35, -27, 12, -28, -14, 8, -26, -45, -31, 14, 5, -6, -21, -6, 5, 11, -4, 45, 3, 21, 8, -28, 33, -4, -3, -14, 5, -12, -11, 14, -25, -43, -1, -22, 14, 12, -29, -24, 12, 8, -6, 20, -3, 4, -25, -1, 10, -1, -8, 7, -3, -15, -19, -26, 20, 15, -30, 30, -4, 7, 13, -3, -20, 11, 23, 20, -1, 27, -24, -14, 11, 7, -35, 31, 10, -45, -42, -8, 12, -3, -13, 48, -3, 22, 5, 2, -20, 12, -7, 25, 13, 19, 0, 8, -2, 10, -15, 12, 15, -36, -35, -6, 16, -14, -4, -6, 13, -17, -15, 10, 4, 3, -4, 4, 12, 12, -1),
    (-9, 10, -16, -13, -14, -4, -4, 21, 1, -28, 4, 27, -4, -6, -6, 7, 5, 15, -19, -13, 12, -4, -36, -12, 4, 13, 12, -42, -15, -13, 13, -3, 4, 27, 0, 41, -9, -3, 34, -5, 7, 8, 7, -14, 11, -3, -33, 13, 3, -4, 19, -29, -9, -4, 20, -17, 2, 30, -10, 31, -15, -4, 21, -17, 4, 12, -12, 9, -4, -1, -35, 22, -34, 21, 2, -35, 4, 10, 14, 9, -4, -9, 11, 20, 13, 13, -27, 36, 15, -1, -20, 3, -7, 23, -6, -34, -28, 20, -1, -51, 8, 14, 11, 20, -20, -30, 16, 33, -3, 4, -11, 37, -1, 12, -26, 0, -31, 32, 5, -24, -27, 12, -10, -45, 11, 4, 12, 6, -20, -38, 19, 28, -18, -20, -17, -5, -14, -1, -20, 1, -28, 16, 19, -10, 2, -5, -3, -7, 11, 12, -31, -4, -10, -9, -4, -25, 32, 42, -56, 30, 1, -32, 6, -24, 28, -1, -12, 13, -9, 5, -31, -14, -13, 26, -25, -15, -18, -6, -4, -25, 7, 36, -5, 8, 1, -8, -14, -3, 4, -3, 10, -9, -20, 22, -19, -17, -11, 14, -13, -3, 8, -1, 12, -2, 4, 12, 9, -4, 7, 1, -23, 1, -17, -12, 2, -51, -8),
    (-11, 14, 30, -11, 22, 4, 27, -12, -11, -6, -9, -15, -11, 2, -14, -4, 0, 15, 16, 20, -29, 14, 21, -4, 3, 10, 29, -5, 34, 14, -4, 1, -1, -1, -15, -11, 14, -4, -44, 21, -8, 8, 36, 20, -27, 4, 31, -4, 13, -2, 3, 4, 18, 17, -9, 4, 32, -13, 7, -13, 23, -5, -27, 30, -9, -10, 17, 4, -28, -12, 27, -10, 15, -5, 19, 4, 12, 23, 4, -4, 13, -13, -25, -44, 16, 14, -23, 1, -16, -5, 29, 18, -23, 9, 29, 8, 25, -5, 7, 21, 34, 14, -29, 18, 28, -17, -32, -56, 17, 13, -60, 3, -12, -32, 5, 25, -12, -5, 6, -8, 23, 2, 8, 14, 12, -20, -28, 28, -38, -1, -10, -29, -4, 7, -12, -3, -18, -18, -6, -19, 17, -26, -18, 8, 20, -14, -34, 3, -8, -9, -34, 18, -4, -4, -5, -15, 7, 4, 7, -4, -15, -8, -22, -29, 6, -15, -4, -2, 14, 0, -7, -16, -30, -1, -24, 33, -4, -26, -9, 19, -18, 1, 4, -2, 1, 12, -45, -5, 5, -13, -20, -22, -57, -17, -19, -13, 5, -14, -20, 30, -37, -40, -7, -3, 17, 12, 6, 14, -21, -26, 22, -12, -9, 0, -17, -8, 1),
    (-17, -14, 19, -5, -9, -32, 2, 2, 12, -38, -18, 16, 3, 11, -45, -2, 20, -21, 1, 21, 28, 6, -5, 28, -37, -14, 34, 5, -4, -46, -7, 4, 4, -62, 4, -7, 8, 23, -13, 10, 9, -7, -4, 5, 30, -12, 14, 41, -33, -16, -2, -6, -26, -39, -34, -7, -14, -37, 20, -13, -11, 9, -15, -6, -16, -19, -6, -6, 0, -5, 18, -3, -19, -21, 23, 23, 20, -19, 15, 0, 1, 0, -13, 25, -9, 3, -4, -8, 4, -10, 1, 5, 5, -5, -5, 37, -14, -25, 50, 27, 36, -25, 11, 6, -14, 6, 11, 28, -30, 8, -6, -33, 23, -11, -20, -10, 24, 7, 2, 59, -11, -25, 31, 17, 17, -4, 4, -2, -4, 9, -8, 8, -3, 3, 12, -27, -27, 15, -21, -36, -22, -5, 7, 44, -23, -3, 3, 22, -4, -9, 9, 7, 12, -12, 11, 21, -11, 12, 5, -2, -11, -20, 4, -7, -3, 12, 10, 22, -8, 2, -13, 16, 18, -21, 12, -5, -13, -5, 10, 26, 5, 14, -10, -19, -24, -17, -19, -15, -9, 15, 4, 27, -7, -35, -22, 22, 21, -6, -10, -14, -10, -13, 11, 18, -30, 34, -12, -5, 3, -13, -30, -45, -35, 5, -7, -16, -2),
    (-6, -12, 11, -1, -31, 27, 11, 0, -35, -4, 26, -1, 12, 19, 19, 17, 14, -20, 19, 9, -3, 19, 9, -11, -17, 17, 9, -19, -39, 17, 27, 0, -29, 10, 45, 14, 33, -7, 57, 20, 21, 13, 21, -5, 8, 2, -11, -35, 11, 23, -10, -40, -38, -1, 13, -9, -24, 15, -2, 10, 2, -29, 14, 15, 9, 8, -2, -22, -10, -30, -12, -46, -22, -29, 10, 13, -27, -3, -29, -15, -8, -33, -5, 13, 33, 59, 8, 20, 9, -27, 25, 3, 5, -17, 5, 11, 3, -23, 23, 7, -41, 3, -11, -21, -5, -39, -2, 18, 13, 28, -1, 18, 3, -18, 21, -7, 34, 0, -12, 31, 4, -28, 11, -5, -60, -7, 1, -3, -3, -39, -29, -3, 5, -18, -25, -12, 3, -4, 14, -2, 6, 11, -30, 12, 1, -17, -16, 3, 2, -6, 4, -5, 15, 10, 13, 6, -14, -16, -29, -36, 27, -4, -1, -20, -20, -36, -31, 0, 5, -11, 5, 8, -10, 3, 19, -4, 21, 15, -13, 35, -15, -19, 6, -1, 28, 23, -14, -2, -5, -1, -30, 28, 3, 8, 6, 9, 14, -6, 38, -10, 13, 3, 3, 31, -11, 7, 0, 0, 5, 7, 5, -15, -14, -6, -12, 35, 17),
    (9, 7, 2, -50, -6, -22, -35, -36, 0, 36, 19, 29, 8, 36, 1, -11, -1, -22, -12, -33, 7, -10, -19, -24, -6, 13, -30, 20, 5, -27, -4, -29, -16, -10, 21, -18, -4, 0, -43, -22, 2, -5, -43, 25, -23, -6, 18, 10, -12, 26, -33, -1, -2, 4, 11, 0, -11, -8, 21, -19, 6, -19, 11, -27, -6, 21, -21, 13, -13, -16, 2, 0, 8, 2, -21, -36, -4, -3, -11, 9, -42, -48, 37, -24, 22, -3, 5, -3, 20, 4, -16, 3, 9, 2, -17, -8, -7, 25, -15, 17, 9, -38, 22, -4, -34, -20, 35, -23, 6, -51, -16, -36, 1, 7, -4, 4, -19, -24, 3, -14, -13, 17, -16, -3, 0, -34, 4, 7, -15, -16, 44, -5, -7, -42, 8, -24, -8, 21, -7, 11, -27, -25, 6, -18, -10, -2, 17, 0, -5, -3, -1, 6, -21, -40, 13, -4, 2, 11, 1, -10, 4, -6, -3, 23, -18, 2, -9, 1, -4, 20, 17, 12, 5, -19, 18, -9, -20, -3, 10, 2, 2, -12, 21, -13, 0, 25, 7, 6, -10, -1, 3, -28, -13, -1, 2, -2, 6, -20, -5, 2, -2, -23, 22, 4, 2, -29, 23, -24, 2, 9, -4, -9, 10, 8, 10, -16, 5),
    (12, -16, -15, 15, -5, -1, -3, -18, 2, 20, -17, -3, -24, 0, 16, -16, 17, -13, -1, -6, 13, 6, -20, 20, 28, -13, -9, -5, -12, -12, 13, -16, 29, 16, -24, 4, -40, -17, -4, -14, 30, 20, 7, -10, 5, 25, -13, 34, 15, 4, -13, -26, 4, -12, -3, -9, 12, 4, -17, 36, -16, -35, -29, -16, 19, 15, -1, 2, 4, 28, -23, 36, 15, -11, -1, -39, -4, -21, 27, -38, -4, 18, -24, 35, -29, -38, 10, -23, 18, 0, 17, -9, -14, -1, -25, 13, 16, -16, 23, -36, 21, 0, 32, -13, 24, 23, -21, 36, -29, -45, -27, -5, 19, 18, 37, -29, 3, 13, -5, 15, 0, -12, 19, -29, 21, 3, 18, 15, 14, 20, -20, 21, -17, -29, -23, 8, 18, 6, 25, -7, 1, 15, -7, 28, 3, 10, 26, -12, 18, 16, 12, 9, 5, 19, -7, 20, 8, -26, -1, 17, 7, 20, 6, 4, -19, 5, -5, -12, 2, -4, 6, -13, 29, 12, 6, 26, 20, 20, -9, 9, -2, -17, -20, 21, 27, -2, 35, 1, 3, 12, -5, -11, 29, -17, 13, 4, 20, -3, -3, 27, 5, 20, -7, -27, -10, 4, -18, 11, 8, -5, 23, 6, 4, -1, 4, -6, -3)
  );
  ----------------
  CONSTANT Layer_6_Columns    : NATURAL := 4;
  CONSTANT Layer_6_Rows       : NATURAL := 4;
  CONSTANT Layer_6_Strides    : NATURAL := 2;
  CONSTANT Layer_6_Activation : Activation_T := relu;
  CONSTANT Layer_6_Padding    : Padding_T := same;
  CONSTANT Layer_6_Values     : NATURAL := 32;
  CONSTANT Layer_6_Filter_X   : NATURAL := 3;
  CONSTANT Layer_6_Filter_Y   : NATURAL := 3;
  CONSTANT Layer_6_Filters    : NATURAL := 32;
  CONSTANT Layer_6_Inputs     : NATURAL := 289;
  CONSTANT Layer_6_Out_Offset : INTEGER := 6;
  CONSTANT Layer_6_Offset     : INTEGER := -1;
  CONSTANT Layer_6 : CNN_Weights_T(0 to Layer_6_Filters-1, 0 to Layer_6_Inputs-1) :=
  (
    (-63, 26, -60, -26, -44, 9, 49, -51, -21, -29, 22, -4, 0, 36, -30, -17, -14, -37, -26, 11, -52, -33, -39, 64, 5, -3, -27, 9, 14, -43, -28, -35, -94, -2, 36, -15, 7, -62, -43, -36, -38, -37, 47, -8, 40, -7, 12, 17, 56, 41, -6, 22, -53, -40, -1, 24, -47, 28, -11, 44, 5, -76, -39, -23, -81, -10, 41, 15, 7, -37, 26, -37, 9, -32, 7, 10, -35, 25, 24, -44, -88, -10, -17, 20, 8, -15, 19, -18, -6, -6, -27, -11, 3, -37, 22, 21, 5, 10, -42, -2, -5, 28, -13, -15, -55, -41, 33, 16, 0, -14, 45, 13, 4, -26, 8, 1, 24, 9, -73, 16, 44, -21, -73, 23, -34, 30, -21, -11, -9, 12, -46, -23, -35, -2, 51, -52, 21, -76, 11, 12, -20, -8, 106, 18, 11, -43, 17, 35, 17, 65, -5, 42, 18, -39, -54, -41, -3, 36, 6, -19, 7, 38, -10, -29, -93, 1, 36, -11, 20, -3, -59, 39, -20, 12, 48, 4, -10, -8, 6, 20, -9, 4, 18, -9, -26, 38, 28, -60, 16, 22, -8, 31, -9, -15, 15, -5, -9, -41, 8, -57, -7, 7, -4, 28, 36, -19, 5, -13, 51, -56, 29, -27, -11, 44, 0, 7, 8, -33, -3, 8, -24, 10, 34, 41, -25, 1, -22, 9, 5, -43, -4, 7, 10, 15, -24, 46, -41, -25, -32, -12, 40, -28, 30, -10, 25, 19, 41, -5, -26, -1, 41, 16, -33, 22, 12, 57, -15, -27, 23, -40, 39, 77, -36, 8, -1, -3, 20, -26, 26, -20, -67, 19, 7, 5, -19, 24, -18, 17, 17, 14, -8, -25, 30, 47, -4, 20, -57, 85, 9),
    (-11, 7, 34, 49, -11, 42, 36, 5, -6, -5, 13, -21, -43, -14, -11, 10, 37, -39, 38, 52, -6, 25, 16, -17, 17, 41, -5, 13, -16, -30, 4, -38, 13, 6, 44, 72, -67, 63, -2, 4, -4, 9, 26, -6, -43, 3, 1, 9, 51, -58, -27, 41, 10, 17, -73, -34, 34, 40, 13, 9, -8, -50, 7, -12, 1, 35, 21, 33, -26, 25, 15, -51, 15, 38, -21, 5, -12, 28, -23, -24, 20, -13, -61, 31, 15, -26, -56, -1, 32, 35, -21, 23, -5, -49, 7, 9, 25, 8, -12, 36, -13, 54, -5, 2, -25, -48, -37, 10, 30, 24, 14, -22, 27, 6, 17, -68, -33, -9, -68, 36, 18, -36, -28, 11, -26, -77, -8, -75, 14, -5, -4, 53, -51, 75, -28, 15, -3, -43, -56, -40, 72, 15, 0, -57, 30, -34, -21, -41, 19, -22, -43, -22, 13, -11, 13, 38, -47, -68, 38, -65, 7, -8, 11, 30, -58, 15, -36, 11, 11, -29, -2, -28, 7, -5, -24, -62, -30, 44, -72, 8, 33, -38, -24, 11, 53, -20, 14, 48, -54, -29, 21, -8, 12, -20, 39, 2, 35, -44, 25, 56, -13, -5, 0, 25, 21, 26, 5, -7, 18, 57, 3, -58, -30, 8, -45, 28, 8, -5, -50, 27, -22, 10, -8, 13, -1, -5, -9, 8, -10, -20, -7, 48, 16, -12, -17, 38, 31, 35, 64, -72, -6, 45, 17, -27, -9, -2, 6, 54, -27, 19, -26, 44, -31, -3, 9, 12, -24, 23, -43, 15, -22, 7, 22, 67, -16, 8, 40, 62, 15, -21, 23, -34, -23, 8, -25, -14, 77, -22, 19, 21, -73, -14, 8, -5, -26, 14, -83, 23, -14),
    (-24, -16, -7, 0, 9, -40, -19, -15, 31, 19, -5, 55, -5, -31, -24, -50, -19, 95, -9, 38, -25, -44, -38, -45, 22, 12, -59, 2, -34, 4, -11, -38, -9, 0, 57, 28, -4, -4, 29, -41, -33, 24, 10, 21, 37, -21, -25, -49, 17, -19, 16, 48, 9, 0, 2, 29, 42, -11, -37, 24, -65, -9, -25, -47, -34, 21, 48, 35, -11, -2, 61, -26, -50, -5, 8, -22, -4, -67, 5, -25, 9, 4, 60, 33, 33, 17, -14, -13, 22, -21, -9, -21, -43, -50, -31, -22, 6, 1, 56, 36, 31, 34, 1, -34, 1, -8, 30, 9, 20, -30, 62, 8, -29, -58, 39, 44, 8, 40, -40, 37, -9, 8, -32, -58, -31, -23, -8, -23, 8, 27, 56, 71, 29, 55, 6, -30, -8, 5, 84, 1, 14, -51, 40, -40, 18, 27, 54, 67, 55, 63, -24, 42, -13, 30, -33, -6, 6, 3, 15, 5, 1, 50, 54, 26, -17, 60, 33, 9, 9, -25, 33, 15, -6, -45, 20, -30, 54, -7, 62, 27, 56, 69, 22, -1, 14, 11, 6, -18, -16, 13, 21, 10, 28, 30, -20, -34, 23, -11, 11, 21, 10, 23, 9, 26, -5, -10, 9, -56, 32, -17, 36, -29, -8, -30, 10, -31, 19, 17, 17, -1, -5, 3, 3, 22, 23, 51, -28, -35, 69, -9, -42, 40, 12, 5, 42, -5, -5, -24, 29, -57, 13, 14, 18, -23, -66, 5, -7, -8, 6, -61, 6, -24, 8, 7, -2, -43, 11, 40, -96, -17, 33, -27, 2, -14, -46, -4, 8, 15, 33, -16, -14, -26, 25, 40, 11, -7, -22, 13, -1, -10, 15, 32, -17, -9, 25, -32, 22, -51, -10),
    (-13, 27, 36, 2, -7, -1, -23, 10, 29, 42, 23, -12, -32, 43, 1, 45, 28, 4, -26, -13, -53, -38, -17, 8, -14, 45, 33, -61, 39, -51, 62, -9, 10, 38, 22, 36, 34, 11, -23, 35, 7, 40, 45, -11, 41, -16, 55, -33, -6, 7, 1, 14, 24, -26, -14, 15, -27, 6, -49, -69, -20, -32, 28, -42, -64, 26, 33, 7, 22, 27, 12, 8, -5, 31, 7, 10, -22, -4, 12, -37, -31, 28, -69, 32, 38, -11, 31, 36, -56, -36, -10, 8, -7, -52, -21, -37, -16, 52, -52, -41, -66, 13, 43, 73, -9, -1, 22, -34, -6, 76, -3, 8, 1, 4, -58, -88, -22, -28, -10, -8, 39, 28, 26, -74, -21, -9, 21, -37, 25, 40, -6, -1, -76, -12, -32, 12, 18, 5, -45, -23, 22, 44, 35, 7, 24, -28, -40, -43, -9, -9, -64, -8, 68, 4, -4, -59, 1, -60, 13, -42, 17, 29, -49, -9, 8, -17, 41, 12, 8, -12, -11, -5, 61, 27, 30, -17, 2, -3, 25, -7, 37, 61, -15, -20, 17, 17, -33, -25, -35, -34, -17, -7, -3, -25, -17, -37, -7, -8, 43, 12, -4, 0, 10, -48, 21, 19, -9, 6, -19, 17, 3, -35, 34, 9, -5, -41, 1, -25, -24, -29, -10, 31, -22, 25, -9, -27, -49, -50, -8, -50, -3, 33, 20, -4, 11, 21, 18, 2, -43, -22, 44, 36, -31, -40, -19, 14, 51, -12, 35, -17, 43, -22, -55, 13, -18, 7, 15, -39, 10, -58, 8, -12, 26, 13, 34, 4, 43, 27, 18, -93, -45, -35, 19, 15, 74, 1, 16, -16, 39, -30, 4, -12, 60, 5, -8, 3, -48, 5, -18),
    (30, -19, 32, -13, 39, -25, -6, -51, 30, 40, -3, -21, -3, -71, 0, -41, -13, 22, 54, 21, 22, 7, 26, 20, -33, -14, 58, -2, -22, -18, -41, 21, 20, 23, 18, -15, 63, -8, 39, -50, -4, 89, 6, -4, -48, -44, -8, -47, -39, 6, 59, 14, 2, -2, 7, 11, -31, 19, 40, -9, 32, -11, -44, 22, 42, 10, -7, -18, 23, 5, 37, -66, -6, 85, 6, 20, -28, -10, -6, -6, -17, -15, 1, 7, -11, -8, 7, -25, -52, 12, -30, -24, 17, 6, -53, 23, 56, 68, 52, -1, 23, -11, 12, -31, -34, 108, -16, 8, -49, -37, -6, 8, -31, -22, 26, 46, -4, -13, -36, -61, -18, 55, 41, -7, 23, 13, -74, -39, 20, 39, 65, 31, 7, 24, -19, -34, -88, 89, -15, 56, -22, -19, -1, -36, -1, -94, 18, 57, 8, -24, -15, -48, 10, 71, 41, -7, 39, 56, -65, -17, -2, -27, 7, 5, -5, 51, -9, -19, -15, 40, 25, 11, -8, -17, -16, 26, 22, -8, 30, 45, -2, -35, -23, -8, 23, 38, 18, 7, 10, 8, -26, -7, -44, 11, -28, -35, -17, 11, -11, 28, 11, -24, 31, -22, 3, -26, -32, 17, 5, 7, -50, -25, 8, -18, 16, -35, 8, 14, -12, 9, -12, 38, -5, -23, -16, 5, -6, -40, -38, 24, -38, 12, 59, -18, 38, -29, 9, -14, -43, -15, 7, 16, -37, -16, -1, -25, 6, -41, 18, -3, -15, 47, -22, 6, -24, -22, -5, -26, 16, -12, -20, -5, 57, 25, -18, 3, -7, -8, 30, -20, -5, -6, -12, 10, -40, 21, -21, -50, -36, -27, 10, -21, -4, 26, 5, 29, -71, -41, -24),
    (11, -14, -29, 28, 46, -31, -1, -59, 3, -42, -36, -44, -7, -26, 28, 13, 5, 15, -13, -6, -46, 10, 6, 25, 13, 5, 38, 38, -20, -28, -46, -24, -48, -9, 6, -16, 56, 12, 16, -40, 28, -15, -10, -20, 43, -55, 103, -25, -43, -26, 7, -20, 31, 17, -8, 50, -48, -29, 21, 33, 0, -7, -41, -35, -55, 24, -3, -7, 2, -10, 44, 10, -14, -70, 35, 12, 27, -38, 69, -13, -62, 7, 8, 28, 58, 71, 15, -37, 17, -51, -31, -30, 8, -43, -35, -23, -2, -34, -42, 47, -19, -33, -9, -4, 17, 13, -29, -2, -40, 9, 0, 48, 7, -23, -56, -31, 1, 5, -1, -46, -1, 22, 50, -8, -51, 11, 16, 7, -45, -40, 34, 27, 16, -48, -16, 31, 24, 29, -73, 12, -60, 51, 31, 8, -43, 45, -11, -39, -9, -33, 17, 2, -47, 23, 73, 10, -6, -9, 8, 16, -21, -18, -14, -39, 74, -6, 5, 81, -18, 15, 33, 18, 16, -29, -23, -43, 23, 75, -40, -49, -76, -75, -38, -50, -16, 22, 4, -22, 40, 42, -28, 48, 10, 38, -10, -6, -50, -8, -58, 38, -44, -46, -16, -16, -13, 49, -4, 16, -16, 47, -24, -23, -44, 9, -15, -15, 24, 14, 3, -9, -12, -19, -37, -8, -4, 21, 88, 34, -43, 41, -54, 1, 14, 27, 17, -26, -44, 1, -3, 34, -31, 22, -15, 19, 32, -40, -36, 9, 31, 30, 7, 55, -25, -48, -39, -21, -13, -11, 54, 25, 25, 16, 43, 12, 40, 3, 12, 1, 6, 2, -3, -19, -12, 15, -77, 20, -7, -59, -24, -10, 32, 16, -2, 35, 26, 21, -55, -12, -4),
    (-1, 8, -10, -7, -48, 36, 42, -2, 7, -9, 38, 42, -7, 5, 39, 24, 17, -54, -30, 55, -6, 42, -3, -19, 6, -20, -20, -14, -2, 1, -2, -12, 3, 0, 8, -26, -25, 27, 9, 23, -15, -8, 50, 72, -33, -21, 12, 30, 101, -56, -13, 39, 6, 49, -6, 9, 24, -23, 32, -41, 46, 8, 5, -7, 46, 38, -29, 0, 1, -12, -3, -1, -1, -33, 33, 14, -20, 2, -17, 35, 62, -25, -13, 7, -13, 71, 10, 5, -26, 1, -74, -86, 23, -36, 29, -29, -39, -11, 0, -24, -36, 40, -53, -7, -3, 29, 35, -34, -24, 24, -8, -14, 27, -27, -25, 4, -2, 35, -21, -9, -11, -44, 47, -25, -36, -9, 22, 24, -4, 33, -4, -57, -56, 68, 52, 38, 0, 17, 14, 43, -27, 29, -12, 24, 45, -4, -28, -63, -49, 38, -27, -38, -7, -57, 56, -67, 36, -34, 6, 21, -18, -6, -62, -43, -25, 23, 40, -1, 15, 21, -7, -2, 55, -42, -61, -13, 26, -13, -18, -37, -53, -8, -23, -19, 4, 24, 7, -54, -8, -7, 6, 20, -28, 23, -27, -44, 4, -44, 27, 30, 14, 25, -27, 22, -3, -2, -9, 8, -9, 45, 8, -28, 3, 7, 7, -7, 31, -35, 15, -41, -20, 23, -18, 23, -80, 8, -36, -28, 22, -17, 20, 39, -10, 25, -4, -2, 8, 10, -21, -14, 19, -15, -13, -38, -63, 24, 4, -47, 13, -2, 29, -1, -24, 28, -3, 70, -21, -26, -6, -42, 38, -14, 25, 31, 29, -27, -35, -30, 21, -49, 23, -29, -1, 35, 37, 15, 29, 0, 11, -36, 0, -13, 8, 27, -28, -23, -21, 56, -25),
    (-28, 42, -90, 29, -37, 45, 11, 73, -5, 27, 3, 3, -3, 29, 8, 11, 39, -21, -57, -14, -24, -4, 1, -111, 17, -3, 7, -45, 40, 0, 8, 7, 6, 59, 0, 24, -69, 6, 25, -1, 40, 15, 34, -2, 31, 24, 23, 40, 50, -55, -61, -27, 23, -9, -48, -32, 29, -26, 6, -56, -15, -37, 9, -24, -4, -18, 23, 28, -74, 1, 17, -2, 11, 8, 15, 12, 15, 7, -12, 1, 46, -8, -15, 18, 33, 1, -37, 17, 40, -33, -14, -18, -12, -47, -1, -25, -15, -57, -28, -17, 14, 12, 70, 25, 12, 3, 19, -69, 64, 22, 5, -53, -3, -23, 27, -42, 26, 13, -1, -27, 7, 17, -10, 2, -44, -10, 24, 16, -53, -3, 21, -42, -58, 48, -9, 39, 46, -39, 7, -49, 55, 22, 33, -56, 23, -4, 23, -108, 41, 23, 14, 55, -6, 16, -10, -23, -115, 14, 65, 8, -13, -13, 68, -13, -65, 23, -27, 49, 55, -25, 8, -23, 62, 12, 0, -39, 24, 18, 41, -39, 39, 31, 12, -10, -8, -36, -8, -16, -41, -46, 16, 0, -38, 39, 5, -24, -25, -32, 23, 23, -37, 8, 1, 16, 14, 24, 10, 14, -9, 9, 27, -2, 10, -9, -6, 44, -25, 7, 20, -34, 24, 9, 7, 10, -26, 40, -26, -82, -14, -47, 36, -3, -16, 2, 65, 30, 7, 50, 24, -33, 6, -19, 2, -15, -22, 29, -24, 2, -22, -40, -44, -73, -10, -1, 23, -10, -20, 15, -53, -30, 87, -20, 44, -20, 8, 7, -10, -16, 55, -11, 22, -15, 14, 13, 38, -43, -24, 15, -24, -37, 2, 26, -13, 10, -5, 5, -18, -43, -40),
    (-81, -50, 2, -16, -55, 8, 12, 46, -60, -60, -39, 41, 12, 6, 46, -1, -27, -9, -43, -29, 59, 14, 48, 45, 26, -36, -24, -14, -24, 7, -17, 69, -30, -72, -79, -24, -40, 41, 47, 33, -59, -66, -52, 24, -21, 3, 1, 23, 44, -44, -38, -52, 21, 12, 13, -71, 7, -37, -8, -25, -5, 5, -19, 47, 11, 20, -18, 2, -25, 16, 11, -7, 6, -10, -36, 44, 38, 20, -9, 14, 36, -21, -34, -34, -13, -24, 14, -27, 16, 2, 12, -29, 9, 31, -25, 25, -33, 8, -61, -2, -49, -2, -2, 2, -57, -56, 20, 44, -23, 24, 19, 17, 25, 2, -40, -20, -34, 12, -13, 5, -3, 2, 9, 22, -32, -7, -6, 33, -30, 18, -55, 24, -53, 38, 48, 15, -93, -26, 21, -15, -33, 29, -1, -5, 6, -50, -38, 29, 32, 34, 24, 39, 22, 9, 10, 85, -48, 30, -24, 36, 5, -4, -9, 25, -4, 67, 36, 44, -8, -11, 37, -9, 9, 44, -22, 5, 15, -2, -89, -4, 22, -24, 10, -7, 18, 6, 14, 17, -33, 30, -1, -10, -8, -26, -31, 13, -55, -32, -13, -14, 55, -20, 10, -31, 23, 0, -15, -20, 19, 30, -10, 40, -21, 24, 9, -6, -24, 55, 31, 40, -12, -16, -3, 36, -25, 12, -14, 1, -11, -13, -9, -17, -19, 13, 43, -7, 13, -37, -9, -34, -7, 25, 4, -8, -27, 32, 21, 5, 25, -2, -8, 47, -4, -18, -50, 17, 41, 6, -11, 3, 2, -1, 6, -2, -40, 15, 12, 22, 68, -16, -6, -19, 52, 11, -34, 35, 34, 23, 24, -4, 13, 8, 4, 7, 2, 9, -11, 10, -19),
    (-17, 8, -6, -7, -29, 36, 78, -37, -78, -11, -5, 32, 2, 29, -70, 43, 36, -52, 40, 3, -2, 29, -55, -8, -5, -66, -70, 9, -25, -8, 35, -60, -46, 9, -15, 6, -54, 47, 77, -24, -78, -1, -25, 74, 27, 28, -75, 27, 17, -90, 39, -14, 7, -3, -39, 23, -69, -61, -52, -41, -5, -24, 38, -16, 4, 24, -19, -6, 24, 40, 3, -40, 9, 48, 13, 51, -28, 11, -41, 8, 18, -53, 58, -18, -12, -26, -1, 31, -50, 11, -27, -24, 12, 7, 30, -27, 16, -27, 32, 32, 25, 14, -54, -18, -85, -24, -25, 11, 19, 18, -24, -13, 12, -40, -1, -57, -20, 23, -46, 40, -13, -98, -25, -3, -45, 8, 8, -8, 33, -39, -25, -23, -21, 56, -7, -16, -82, -8, -8, 54, 16, 24, -26, -1, 25, -81, 21, -41, -36, 23, -8, 0, -21, -38, -24, 1, 2, -11, 50, 2, -40, 7, -23, -14, 22, 39, -9, -24, 13, 2, 37, -11, 41, -99, -21, 4, 24, -11, 22, -42, -37, -13, 3, 18, -66, 10, -29, -8, -9, -36, -15, 13, 12, -21, 5, -28, 17, -3, -57, -5, -5, -33, -36, -13, 27, 9, 22, 16, 68, 14, -23, -8, -16, 41, 4, 70, -5, -28, 21, 44, -31, 11, -28, 44, 24, -8, -21, -13, 47, 6, -51, -15, -60, -25, -4, -5, -10, -8, -3, 18, 15, 27, -24, 8, 5, 29, 5, 2, -6, -36, -5, 27, 15, 8, -13, 27, -12, 44, -2, -19, 2, -1, -1, 38, -37, -11, -3, 24, -33, 1, 6, -17, 9, 11, -26, 64, 2, 2, 20, -3, -43, -2, -24, 14, -2, 35, -113, -16, 4),
    (8, -57, -37, 22, -9, -28, -3, 39, 27, 12, -27, -14, -40, 35, -49, -6, -15, -41, -48, -23, 8, -24, -35, -28, -43, 23, -5, -21, -14, 39, 10, 25, -48, -42, -6, 16, 6, -28, -3, 22, 79, -41, -78, -39, -73, 27, -25, -1, -26, 27, -50, -76, -29, -30, 28, -30, 31, 52, 51, 44, 35, 87, 11, 55, -53, -49, 24, -67, 23, -9, 33, 20, 43, 31, -23, -31, -38, -16, -12, -8, -3, 15, -5, -36, -19, -27, 6, -47, -39, 46, 16, 16, 40, 21, 1, 46, 39, -7, 34, 38, -6, 34, -49, -4, 50, -20, -3, -8, 1, -14, -8, -4, -35, -9, -56, 29, -29, -24, 12, 8, 31, 54, 16, 40, -41, -33, -25, 0, 25, -20, 36, 83, 0, -10, -54, -60, 71, -27, -42, -49, -85, -5, 7, -1, 0, 11, -25, 101, 10, -61, -12, 5, 36, 17, 39, 60, -6, -30, -8, 8, 33, -32, 36, 8, -2, -22, -27, -7, 0, -17, -30, 7, 2, -1, 31, -50, -2, -8, -103, 21, 19, -24, -2, 23, 12, -29, -40, 12, -12, -44, 25, -32, 14, 34, -51, 24, -28, 26, -4, -24, -22, -20, 43, 14, 0, -17, 25, -53, 30, 15, -14, -2, -40, -31, -30, 3, 39, 6, -52, -11, 11, -37, 7, -50, 28, 8, -12, 11, -18, -27, 21, -6, 5, -26, 12, 8, 38, -11, -10, -36, -25, 6, -10, -21, 2, -32, -28, -2, 6, -39, -54, -37, -7, -41, -14, -61, -1, 22, -97, -21, -17, 8, -10, -8, -71, -19, 2, 40, 1, 45, 24, -40, -28, 12, -28, -13, -3, 41, -9, 32, -43, 1, 4, -34, 7, -49, 2, -10, -4),
    (33, -27, -9, 2, 18, -12, -6, -21, 23, -31, 1, -8, 63, 9, -18, -22, 10, 10, 10, -8, -35, 12, -40, -25, -77, -9, -56, -23, 25, 4, -24, 21, 5, 11, -29, -46, 50, 8, 16, -29, -11, -56, 25, 10, 54, -33, -8, -41, -10, -7, 6, -7, -12, 1, -8, 26, -61, -40, -39, -27, 27, 5, -6, 18, 16, 6, -28, -19, 35, 22, 15, -58, -23, -43, 10, 39, -49, -13, -23, 6, 10, -24, -14, 9, 10, 25, -32, 4, -60, -26, -10, -7, 11, -1, 14, 9, 28, -33, -39, -69, 50, -24, -18, -18, 13, 11, 12, -14, 11, -9, 9, -30, -8, 4, 11, 27, -25, 24, 41, -11, -81, -10, -27, 36, 67, 75, -45, 48, 8, -28, -1, -91, 81, -10, -19, 7, -10, -6, 69, 9, 58, -28, -6, 8, -8, 32, 21, 41, 12, -5, 60, 25, -57, -43, -4, 48, 73, 90, -9, 22, 9, -16, -31, -27, 33, 33, -7, 36, -29, -6, 29, 18, 44, -26, -11, -11, 28, 29, 30, 38, 15, 41, 52, -9, -46, -25, -19, 40, 18, 103, 58, -9, -75, 8, -59, -25, -12, -17, -16, 32, 6, -8, 22, -48, 12, -40, -12, -32, 4, 39, 5, 35, 1, 0, 27, -41, -9, -49, -38, -3, 38, 55, -62, 39, -26, -41, -59, -83, 75, -36, 34, 36, 27, -33, 22, -31, 26, -17, -33, -11, -37, 48, -8, 25, 48, -22, 7, -5, -24, -31, -13, 13, 37, 40, -31, -7, 1, -30, -74, -47, 70, -38, 27, 0, -14, -25, -3, -29, 18, -54, -23, -71, 9, 48, -1, 46, -54, 6, -11, -38, -9, 16, 13, 13, -11, 30, 20, -16, 47),
    (8, -2, 20, -5, 14, 5, -20, 34, -6, -25, 1, -8, 5, -8, 22, 5, -11, -1, 24, 1, -10, 22, -20, -15, -16, -16, 3, -14, -62, -33, 34, -3, 22, -15, -13, -8, 23, -22, -42, 22, 29, -6, -23, 23, 20, -10, 11, -15, -16, -7, 6, 8, -18, 8, 8, 24, -11, -10, 14, 8, -32, -26, 40, 28, 27, 19, 25, -38, -21, -23, -51, -25, 39, 4, -5, 18, -35, 16, 26, 3, -12, 0, 3, 30, 3, -18, 42, 23, -15, 9, 4, 18, -29, 17, 8, 20, -21, 1, 5, -36, 21, -51, 24, -10, -43, 27, -58, 24, -6, 18, 23, 9, -92, 13, 39, 26, -25, 15, 40, 72, -54, -54, 27, -37, -57, 26, 23, -24, 7, 55, -8, -40, -11, -73, -41, -29, -44, 39, -4, 38, 7, 4, 9, -36, -60, -63, 48, 14, -71, 59, 60, 75, -84, -33, -14, -88, -15, 31, 32, 17, -23, 46, 12, -32, 4, -42, -23, -23, -11, 53, 26, -10, 35, -42, 28, -24, -47, 0, 48, 9, -46, 52, 43, 32, -57, -8, -43, -41, -25, 62, 3, 0, -42, 23, -2, -27, 11, 2, 52, 20, 40, 34, -6, 21, -13, -3, 5, -5, -30, 6, 39, 26, -9, 21, -14, 27, -42, 22, 17, -19, 25, 76, 6, -16, -17, 38, 3, -63, 65, -29, 34, 89, -34, 64, 31, 33, -59, -14, -27, -46, -21, -32, 44, 31, -6, 37, 52, 9, -50, 23, 36, -28, -10, 89, 17, -34, -24, -37, 35, -62, 58, -10, 40, 23, 43, 12, 38, -25, 44, -107, -36, -48, -37, 19, 8, 16, 9, -30, -11, -50, 8, 57, -11, -2, 44, 32, -39, -39, -12),
    (7, -32, -13, 1, -7, 8, 9, -5, -22, -8, -35, -16, -19, 34, -28, 23, -11, -27, -3, -73, -27, 5, 0, -10, 28, -31, 39, 11, 12, 25, 16, 19, -1, 39, -22, -35, -21, -50, -13, 12, 7, 28, -60, -4, -30, 51, 6, -23, -22, -36, -17, -56, -37, 22, 17, 29, -58, -10, 23, -50, -11, 23, 14, 39, 2, 25, -19, -56, -24, 8, 6, -45, -1, 5, -8, 8, 24, 6, 18, -6, -21, -5, -25, -41, 4, -40, -23, -1, 4, 7, -47, -21, 8, 8, -24, 28, 15, -19, 71, 55, 26, -58, -16, -38, -21, -5, -28, 53, 10, -34, 10, -16, -28, -11, 44, 94, 6, 20, 5, -3, -21, -8, 23, 22, -19, -18, -47, -11, 30, -3, 45, 29, 48, -59, -22, -11, -47, 27, -17, 50, -35, -29, 10, 25, -4, -39, 32, 100, 22, 34, 71, 11, 3, 7, 66, -10, -52, 70, -24, -8, -2, 50, -7, 22, 69, -47, 23, 5, -22, 18, 52, 21, -9, -22, -17, -7, 9, -28, 26, 2, -21, -29, 18, -14, -2, -29, 63, -1, -22, 62, -25, -10, -30, 1, -52, 0, -18, -9, 29, 7, -47, 20, -9, 8, -1, -12, -15, -8, -11, 27, -25, 15, -24, -31, -44, -31, 1, 25, -17, -24, 4, -16, 1, -32, 18, -18, -21, -7, 21, 8, 0, -2, -13, -60, 16, -24, 6, -4, -16, -3, -29, 63, -52, -17, -3, -20, -14, -56, -20, 24, 10, -23, -20, -31, -2, -72, -4, -50, 10, -22, 34, 0, 5, 20, -68, -37, -53, -39, 41, -53, -58, -14, -34, 48, -9, 4, -19, -26, -28, -32, -1, 11, -42, 8, 36, -13, -80, -30, -10),
    (-15, 17, -6, -54, -21, 11, 44, 22, 16, -44, -18, -59, -65, 47, -43, 1, -11, -47, -93, -36, -23, -42, 34, 1, -28, 23, 18, -45, 32, 75, 23, 51, 42, 23, -33, 0, -57, 9, 28, 72, 32, -51, -35, -22, 9, 47, -38, 61, 18, -30, -23, -37, -21, -25, -44, -51, -1, 3, 4, -23, 36, -4, 55, 3, -7, -9, -62, -3, -2, 15, -39, 88, 27, -16, -9, 11, 17, 47, 8, -6, 7, -18, -24, -6, 4, -31, 4, -38, 17, -9, 26, -16, -4, 7, 8, -8, -52, -57, 46, 51, 6, -24, -22, 31, 17, -21, -9, -8, 26, -8, -14, -8, -88, 37, -23, -14, 54, -45, -18, -43, 57, 25, 5, -4, 7, 37, -38, 17, -30, -46, -55, -24, -39, -16, 36, 62, 22, -22, -41, 8, 7, 66, -12, 27, -20, -2, -37, -64, -100, -9, 18, 24, -83, -15, -12, -9, 2, 16, 42, 4, -26, -7, -73, 23, 17, -32, -36, -30, -15, -24, -3, -1, 22, 56, 11, -16, -41, -6, 33, -44, -46, -14, -24, 38, -9, -20, 2, -7, 3, -22, 25, -5, -63, -25, 38, 25, 38, -2, -1, 18, -10, -10, -50, -6, 32, -18, -26, -30, -22, 32, 9, 3, 36, 6, -18, -19, 3, 4, 19, -6, -30, -17, -4, -46, -8, -27, 16, 12, -1, -22, 15, 8, 59, 6, 8, 1, -7, 24, 12, 32, -27, -24, -16, 37, -5, 29, -3, 29, -24, 37, -9, -2, 14, 26, 21, -14, -9, 23, 1, 35, 26, -4, -8, -40, 16, 15, -20, -5, -2, 0, 44, 17, 22, -9, 8, 28, -17, 19, 0, 3, 36, -11, -16, -30, -38, 23, 30, -35, -14),
    (-51, -5, 22, 21, -2, 33, -3, -19, -10, -19, 50, 7, -5, 9, -44, -55, 34, -24, -9, 12, -5, -8, 13, -14, -5, 10, -34, 16, -4, -12, 8, 11, -48, 18, 64, 48, -23, -4, 12, 42, 41, -32, 25, 14, 39, -6, -38, -5, -51, -28, -16, 55, 36, -41, 38, -1, 22, 26, -37, -18, -67, -56, -18, -27, -43, 1, 41, -1, -18, -49, 8, 36, 22, 7, -9, -14, 7, -9, 13, 5, 12, 33, -5, 38, 12, -8, 9, -30, 41, 9, 8, 33, -40, -41, -45, -7, -17, -17, -55, -52, 6, -3, 15, -37, -27, -41, -74, 28, 10, -29, 39, 3, 21, 19, 3, -12, 33, 39, 11, 7, -4, -44, 9, 17, 22, 14, -22, 44, 2, 25, -61, -62, 19, 57, 29, -18, -27, -51, 2, 56, -6, -38, 24, 13, 63, 54, -25, -61, 24, 0, 11, 10, 1, -33, 45, -57, -14, -7, -29, 60, 20, 35, -65, -32, 7, 72, 40, -57, -41, -73, -34, 24, 60, -4, 14, -10, 44, 28, 5, -17, -18, -16, -60, -33, 11, -32, -1, -48, 18, 14, -36, 1, -60, 4, -16, -39, -1, 20, 24, 12, 36, 13, -5, -1, -6, -23, 16, -30, 18, -7, 4, -1, -56, -6, 35, 20, -20, -5, -13, 16, -17, 47, -42, 10, -61, 3, 11, -6, 28, -26, -11, 34, 24, 22, -4, 0, 50, -34, 20, -59, -10, -59, 8, 25, -14, 24, 31, 7, -21, -23, -24, 69, 70, 40, -8, 16, -43, -45, 4, -40, 9, -45, 6, 29, -20, 30, 11, -9, -15, -18, 30, -57, 27, -30, 1, 9, -12, 93, 4, 19, 24, -51, 21, 63, -14, 42, -14, -5, 10),
    (-55, 36, 10, 9, -6, 22, 5, 5, 32, -4, 53, 7, -28, -13, -20, 2, -29, -33, -46, 5, -7, -52, 39, -25, 20, -7, -10, -24, -48, 20, 9, -14, -54, 34, 44, 14, -10, 54, 51, 28, -3, -26, 40, -3, -29, 3, -4, -33, 21, 64, -48, -10, 18, 2, -4, 7, -6, 18, -5, 16, -7, 27, -26, -18, 9, 24, -30, -37, 7, 32, 48, -46, 13, 10, 19, -2, 17, 27, -28, -40, 33, 36, -71, -34, -8, 37, 17, 20, 24, 15, 34, -9, 16, 17, -24, 5, -33, -31, -41, -20, -51, 41, 48, 68, -44, -28, 27, 9, -9, 38, -105, 30, 29, 8, -41, -61, 15, -20, 2, -20, 10, 2, 8, -18, -40, 46, 16, 22, -19, -87, -40, 30, -89, 35, 37, 42, -10, -24, -24, 31, -24, 40, -65, -4, 9, 38, -55, -99, -26, -24, -6, -60, 13, 21, 8, -4, 30, 53, 21, 38, -9, -58, -37, 4, 38, -10, -12, -11, 22, 1, 3, 20, 50, 8, -27, 11, 35, 16, 7, -25, -4, -46, -47, -40, 21, 38, 3, 46, 18, 74, -5, 31, -21, -41, -43, -24, 19, 10, -31, 20, -31, -45, 5, 5, 9, 8, -25, -13, 38, 0, -30, -36, -13, 5, -6, -34, 7, 11, -26, 25, -10, -24, 53, 52, 25, -20, -51, 25, 11, 20, -55, -35, -1, -40, -23, 2, 1, 18, -34, 9, 50, 21, -6, 23, -10, 8, -9, 37, 20, -14, -16, 69, 8, -48, 37, 22, 22, -8, -55, 24, -14, -38, 26, -35, 17, 11, 6, 16, 4, -5, -4, 7, 31, 19, -23, 13, 28, -22, -23, 14, 28, 0, -31, 32, -26, -34, 21, 7, -9),
    (16, 3, -14, 19, 2, 21, 10, 10, -4, -20, 5, 5, 22, -35, -14, 23, 16, -25, 10, -49, 6, 9, -28, -12, 15, -20, -30, 6, 65, 15, -9, 23, 12, -13, -24, -12, -15, 49, 55, 2, -32, -48, -7, 21, -18, -20, -36, 39, 36, -39, 38, -39, 36, 42, -36, -29, 68, -7, -63, 10, 6, -9, 18, 23, -19, 6, 34, -45, -23, 33, 40, 13, -25, -52, -10, 1, 26, 21, -30, -9, 23, 9, 17, -21, 20, 19, -34, 9, 43, 8, -30, 48, 7, 37, -14, 48, 10, -71, -13, 24, 24, -52, -72, -54, -42, -4, -55, -23, 22, -41, -19, -53, -2, 5, 33, 36, -16, 29, 2, 8, -20, -12, 10, 45, 42, -29, 7, 24, 15, -79, 46, 27, 45, -53, -84, -77, -43, -8, -24, 40, 17, -56, -26, -40, 20, 16, 38, 1, 26, 9, 7, 18, 1, -34, 35, 70, 16, -29, -15, 23, 13, -4, -28, 10, -35, -25, -49, -33, -54, -13, 4, 14, -29, -47, -11, -40, 15, 23, 30, -10, 16, -10, 13, 41, 26, 14, 42, 33, 6, -2, -25, 30, -71, 52, -7, -33, 33, -9, 7, -72, -31, 24, 16, 55, 8, -10, 24, -59, -92, -10, 10, 23, 23, -33, -12, 46, -29, 22, -26, 9, -12, 8, 32, -55, 3, 24, 17, 4, 56, 23, 46, -21, -60, 16, -24, -8, 6, -58, -2, -17, -41, 31, 43, 23, -10, -16, 0, 24, -21, -14, -35, -16, -8, -9, -8, -75, 9, 47, 18, 2, 43, -7, -4, -1, -76, 5, 29, 16, 8, -12, 26, 3, -25, 11, -14, 38, -9, 33, 37, 25, -14, -39, -27, -27, 22, 9, 18, -60, -18),
    (29, -7, 65, 8, 27, -53, -50, -88, -16, -1, -45, -64, 23, 23, 14, -28, -22, 24, 27, -2, -67, 6, -11, 1, 16, -3, 14, -2, -4, -35, 10, -63, 30, -6, 7, 36, 39, 1, -20, -29, -80, 17, -44, 29, 41, -14, -58, -23, -4, -73, 26, 23, 20, 17, -29, 46, -11, -11, 16, 29, -38, -32, 67, -66, -14, 23, -37, 32, -54, 11, 1, 12, -54, 1, 20, 28, 9, -10, -27, -2, 6, -48, 32, 12, 54, 9, -5, 15, 5, -41, 31, 28, -64, 3, 19, -9, 3, 10, -38, -15, 6, -24, -47, 47, -27, -28, 23, 5, -24, 30, 11, 15, 36, 53, -30, -19, -32, -6, 7, 44, 17, 16, -27, 37, -37, 23, -11, -20, 56, 18, -7, 0, 56, -30, -62, 19, -21, -55, -34, 1, 23, 48, -4, -35, 35, 3, 10, -40, -78, 14, 5, 24, 22, 16, -43, -5, -41, -53, 31, -34, -19, 44, -13, 39, -3, 46, -16, 5, -5, -47, 32, -22, 37, -16, -31, -37, 2, 19, 5, 51, 29, 36, 4, 8, 57, -16, -74, 3, -30, -37, 66, -57, 26, 6, -15, -36, -18, 32, 17, 23, -12, -26, -52, 11, 1, -11, 43, -105, -17, 60, -28, 24, 33, 15, 9, -16, 9, 34, 39, 41, -4, 32, -62, 13, 18, -14, 12, -57, 33, 32, -44, 35, -29, -18, 31, 37, -30, 40, 19, -24, -2, 5, -3, 5, 15, 14, 62, -9, -33, 30, 42, 28, -29, 42, -31, 27, 38, 24, -48, -10, 30, -1, 21, 45, 2, 5, 22, 22, 38, -38, 3, -86, 10, 16, 4, 25, -28, 13, -19, -16, 15, 15, -27, -12, -38, -43, -58, -6, -1),
    (-11, 17, -2, -7, 20, 36, -14, -19, -6, 51, 17, -15, -22, -51, -37, -11, -24, 3, 23, 36, 5, 29, 30, 28, -29, -41, 24, 19, 5, 54, -18, -8, -24, 58, -20, -16, 15, 73, 54, 20, -11, 27, 44, 37, -24, -25, -6, -10, 10, -24, 24, 64, 32, 11, 20, 15, -25, -30, -28, 13, 52, 71, -28, 6, 15, 5, -7, -36, -13, 40, 49, 6, -3, -28, 24, 16, 7, -7, 16, -13, 1, -12, 1, 23, 37, 24, -7, -12, -18, -7, 16, -5, 26, 22, -15, -1, -45, -4, -14, -25, 13, -30, -7, -45, 20, 60, 0, 2, 34, -39, 5, -29, -4, -1, 30, 32, -33, 15, -4, -3, -8, 8, -10, 3, -26, 17, -8, -23, -51, -42, 20, -67, 40, 30, 48, -37, -47, 43, 91, 43, 29, -86, 7, -47, -9, -39, 26, 29, 48, 39, 23, -28, -9, -48, 30, -10, 24, 66, -41, 10, -37, 38, -15, -82, -10, 70, 45, 59, -18, 33, 48, 24, 17, -76, -8, 7, 31, 17, 77, 0, 6, 73, 25, -21, 9, 6, 26, -23, 23, 45, -51, 35, -30, 9, -63, -50, -29, 10, 19, -44, -48, -38, -6, -37, -21, -28, -7, -25, 36, 9, 6, -12, -9, -21, -60, 6, -7, 9, -39, 12, 27, -24, 14, -11, -59, 28, -71, -17, -7, -8, 62, -4, -25, 24, 29, 65, 23, -37, 44, -9, -54, -7, 40, -1, 36, -24, 7, -24, -2, 1, 22, -37, 21, 22, -20, -19, -36, 2, -1, -48, 7, -21, 24, 47, 19, 8, 37, 52, -5, 0, 2, 10, -8, 33, 27, -9, 15, 12, 24, -44, -7, 13, 28, -23, 32, 24, -68, -29, 17),
    (-9, -9, -53, -36, 25, 17, 8, 56, 39, 8, -13, -10, 1, 9, -43, -9, 16, 47, -40, 1, 14, -4, 20, 34, -2, -5, -33, 50, 17, 10, 8, -5, -46, -4, -43, -50, -35, 7, -8, 35, 45, 2, -22, -78, -22, 42, -13, 30, 20, 23, -38, -2, -7, -28, -47, 0, -19, 9, 1, 61, -2, -24, 25, 36, 8, -19, -12, -7, -4, -14, 14, -16, 57, -1, -34, -22, -35, 56, 20, -67, -77, 17, -78, -8, 21, -6, 36, -7, 28, 2, 39, 11, 26, 22, -11, 0, 22, 8, 44, 11, 76, -13, -70, -24, -1, 2, -22, -23, 24, -73, 17, -33, -43, -82, 16, 5, 11, 24, 51, 55, -31, -71, 3, -5, 39, -2, -23, 20, 8, 8, 25, -56, -11, -9, 5, -5, -25, 66, 13, -17, -33, 6, 21, -1, -23, -55, 38, -7, -6, 8, 30, 40, -104, 23, 32, -48, 14, -17, -15, 34, 11, 56, 4, 9, -15, -25, -13, -55, 13, -38, 11, 23, 34, -11, 9, 6, 14, -57, -64, -41, -53, -28, -45, 9, -27, -14, -9, -82, -3, -49, 22, 27, -59, 29, -33, -15, 10, 8, 24, 32, -57, 56, 32, 16, 36, -21, 12, -59, -55, -43, 47, 16, -10, 1, -58, -43, 22, -43, 35, 5, -34, -13, 8, -40, 22, 26, 28, 13, 27, 25, 39, 29, -11, 51, 28, 14, 15, -51, -11, -40, -36, -47, -16, 72, -1, 21, 16, -21, -20, -53, 4, 1, -6, 84, -39, -54, 20, -7, -12, -7, 5, 12, 34, 39, -2, 21, 27, -10, -13, -72, -63, -16, 46, 11, -8, -16, -46, -9, 45, -24, 1, 16, 79, 31, -18, 11, 24, -6, -4),
    (42, -8, 12, 10, 33, -15, -25, -25, 8, -10, 54, -14, -3, -41, 11, 18, -10, -32, 47, 7, 36, 20, -40, 4, 0, 23, -43, -51, -21, 2, 17, -21, 24, -2, 68, 1, 11, -4, -33, -43, 11, 26, 27, -18, 16, -6, 42, -23, 57, 8, 56, 20, 32, 88, 13, 41, 5, 8, -13, -26, 19, 1, 25, -6, 32, 22, -24, 7, -17, 8, -39, -3, -3, -10, -30, -17, -39, -32, 35, 1, 28, 29, -40, -13, 4, 70, -15, 22, -24, -31, -11, -6, 46, -29, -13, 11, 21, 3, 31, 25, 17, -8, 14, 1, 35, -9, -22, -8, 19, -28, 49, -12, -33, -45, 54, -19, -12, 26, 24, 1, 11, -25, -7, -40, -34, 57, 7, -10, 16, 32, 1, -55, 4, -28, -40, 84, 40, 25, -9, 23, -41, 24, 34, -14, 2, -21, 43, -38, -81, 20, 45, -39, -8, 4, 24, -47, 25, 29, -4, -28, -12, 23, -16, -65, -19, -39, -42, 56, 15, 12, 15, 10, 19, 27, -34, -23, 7, 33, -23, 3, -28, -17, 25, -60, 13, 21, 52, -26, 36, 9, -82, -8, 14, 6, 6, -11, -67, -19, 12, -10, 32, 25, -2, -5, -50, 12, 0, -25, 15, -23, -17, -9, -9, -41, 2, 30, -5, 43, -37, -41, -3, 1, -7, 23, -79, -1, -48, -10, -7, -10, -11, 23, 15, 44, 8, 20, -10, 12, -14, -2, -19, -64, -49, -45, 39, -56, 10, -91, -45, 26, 11, -38, -9, 27, -24, 21, -29, -6, 43, -51, 34, -9, 9, 10, 56, 52, 23, -2, 29, 27, -37, 24, 5, 29, -7, -14, 55, -20, 24, -11, -31, -10, 23, -19, 14, -13, -20, 53, -1),
    (26, -14, -20, -7, -41, 7, 9, 9, 4, 28, 1, -27, 0, 42, 5, -23, 40, 25, -24, -1, -11, -14, -25, -40, 20, 22, 25, -8, -2, 27, -9, -8, 8, -43, -8, -12, -10, 8, -23, 22, 27, -4, 5, -48, 13, 28, -41, -16, 39, 61, -36, 22, -26, -10, -25, -47, 43, 54, 14, 31, 25, -18, -8, -11, 11, -42, -13, 34, 10, 23, 12, -49, 1, -27, 8, -35, 10, 6, 8, -21, 25, 22, 7, 28, 18, -13, -45, 27, -8, 49, -19, 50, 4, 9, 15, 5, -30, 23, -5, -26, -58, 39, 16, 25, 20, -12, 25, -69, -8, -3, 41, -25, 21, 31, -40, -21, 10, -25, 17, -29, 36, 20, -19, 10, 19, 16, -39, 12, -10, 54, 22, -13, -41, 28, 12, 39, 71, 8, -3, -42, -20, 5, -7, 43, 40, 69, -89, 2, 9, -51, -22, -79, 95, 70, 24, -10, 68, -17, -68, -40, 24, 25, 7, 4, -14, 23, 1, -16, 36, -7, -18, 8, 66, 44, 1, -14, 44, 2, -21, -24, 5, -38, -21, -48, 106, 42, 10, -15, 87, -20, -6, -10, -48, 22, -79, -42, -26, 29, 25, 10, -13, 5, 43, 19, -26, -30, -5, -46, 31, 4, -22, 20, 35, -44, -34, -38, -15, 3, -2, 12, 9, 0, -38, -56, -58, 26, -98, 12, -49, 6, 14, 41, -7, 8, 44, 2, 15, 22, -30, 11, 24, 19, -89, -24, 2, -55, -25, -55, -1, 16, -28, -39, 37, -14, -39, -47, -7, 56, -25, -42, -19, 13, 22, -32, 7, -5, 8, -19, 29, 15, -9, 41, 32, 60, 41, -1, 18, -21, -20, 5, 24, -8, 5, -21, 29, -40, 19, -10, 0),
    (-8, -31, -26, -21, 21, -17, -8, 0, -7, 45, -29, 47, 13, -14, -11, -7, -39, -36, 13, -15, -3, 5, 51, -22, -2, -52, -26, -12, -25, 2, 38, -3, -32, -50, -27, -74, -25, 7, -20, 31, -16, 69, 12, 23, 2, -5, -14, 1, -14, -11, 18, -1, 53, 34, 79, 27, -15, -87, -29, -14, -28, 5, -17, 29, -75, -16, 28, -35, -10, 30, -22, -37, 54, 45, 23, -20, 5, -41, -19, -33, -5, 31, -11, 9, 14, -45, 14, -21, -46, -12, 0, -16, -8, 1, -50, 61, 2, -32, -12, 7, 40, -59, -53, 0, -28, 17, -51, -30, 32, 16, 20, 1, -24, -55, 1, -90, -6, -6, -25, 74, -59, -25, -11, 7, -47, -8, 34, 13, -11, -8, -24, 7, 0, -57, -36, -33, -37, -52, -28, 9, 72, 4, 39, 7, -8, -14, 8, -55, 25, 22, -11, 80, -60, -103, -63, 8, -69, 8, 30, 39, -62, -44, 7, -12, 1, 31, 5, 38, 11, -60, 7, 5, 37, 8, -23, 5, -22, 22, 23, 62, 37, -2, 57, -45, -70, -13, -2, 35, -14, 51, -1, 36, 13, -10, 30, 6, 5, 23, -20, 32, -6, 25, 3, 32, -3, 37, 28, 41, 12, -4, -3, -6, 8, 12, 9, 22, -8, 8, 31, 14, -38, 34, 14, 3, 24, -26, -65, -5, 21, -16, -57, 5, 5, -23, -36, 17, 20, 44, 42, -1, 21, 42, -9, -31, -58, 42, 27, 31, 5, -10, -41, -5, -39, -8, 29, 35, -13, -14, -33, -15, 10, -31, 37, -26, -5, -53, 3, 34, 34, -74, 60, -30, -21, 42, 28, -13, -37, 22, -19, 5, -9, 67, -111, 19, -8, -10, -35, -16, 38),
    (-50, 7, -14, 0, 13, 23, 57, 5, -3, 38, 18, 20, -21, 20, 41, -40, 19, 37, -4, 11, 10, 8, -20, 5, 17, 44, -38, -21, -7, 45, -5, -39, 5, 40, -10, 23, -8, 2, 36, -5, -8, 25, 32, -17, -20, -21, -7, -17, 37, 19, -3, 59, -24, 21, 11, -28, 42, 7, -8, -12, 34, 10, -12, -57, 17, 18, -3, 23, 7, -3, 3, 0, -29, -7, 0, -1, -12, -23, 9, -25, 37, 34, 27, 8, -32, 7, -15, 1, 61, 32, -20, 14, 21, 7, -58, -28, -26, -68, 6, -43, 6, -38, -37, 10, -6, -2, -19, -12, -21, 6, 24, -28, -48, -44, -21, -37, 35, -1, 54, 24, -16, -55, 32, 5, -26, 45, -7, 41, -38, -23, -23, -67, 10, -22, -50, 12, 20, -36, -55, 36, -80, 18, 9, -14, -29, -16, -32, 7, -23, -12, -30, -24, -13, -22, 41, 5, 13, 26, -18, 70, -49, 43, 8, -95, 10, -6, 7, -29, 3, 4, -54, -5, 39, 27, -26, -23, -34, 43, 0, -34, -24, -13, -52, -5, -28, 12, 37, -27, 42, 10, -38, 40, 8, 39, 53, 43, 25, 21, 17, 0, -1, 104, -20, 17, -62, -45, 4, 18, -9, -32, -8, 90, 13, 8, 22, -16, 8, 31, 65, 45, -35, 9, -45, 23, 7, 19, 72, 52, 8, 33, 12, 2, -14, 50, -22, 65, -25, 2, -8, -9, 9, -88, 6, 88, 12, 48, 49, -8, 6, -29, 54, 13, 55, 41, -24, 3, -29, -27, 48, 16, -11, -13, -23, 18, 7, 19, 47, 50, -28, 13, 12, 37, -23, -33, -39, 20, 11, -35, 12, -19, 3, -10, 8, -9, 7, 6, -42, 20, -1),
    (35, -10, 28, 15, 22, -33, -52, -21, 76, -5, -14, -60, -6, -26, 19, -70, 17, 71, -22, 4, 10, -45, -21, -21, 22, 33, 9, 40, 23, -7, -9, 63, 24, -60, 40, 14, 36, -6, -19, 41, 93, 8, 6, -60, 9, -33, 55, -60, -46, 69, 2, 38, 28, -53, 39, 19, 3, 13, 16, 26, -65, -60, -75, -13, -51, -44, -6, 17, 22, 10, 8, 9, 6, 18, 9, -31, 26, -19, 65, -45, -4, 7, -60, 10, 31, -24, 22, 5, -17, -47, -46, -2, -52, -16, -40, -34, 5, -13, 41, 29, 19, -1, -42, 21, 81, 20, 0, -90, -5, -12, 6, -38, 9, 32, -38, 42, 20, -41, -6, 5, 20, 26, 12, 35, 6, 52, 16, 38, 9, 17, 28, 9, 67, 11, 19, 21, 60, 11, -11, -26, -5, 1, 0, -36, -7, 29, -8, 24, 40, -8, 5, 1, 26, 60, -7, 22, -60, -6, -8, -5, -7, -36, 33, -11, 38, -12, 57, -24, -4, 11, 60, -29, 56, -4, 8, -26, -12, 82, 43, 36, 20, 9, -13, 15, -24, 7, 6, 10, -56, 2, 24, -17, -5, -23, 55, 3, 4, 18, 64, 14, 19, -21, 15, -61, 34, -23, -3, -33, 7, -47, -36, 4, 19, -11, -2, 3, 31, -4, -24, 22, -10, 16, -39, 21, -16, 10, -13, -25, 16, 24, 33, 1, 48, -25, 15, -8, -7, 19, 6, -41, 14, 6, 6, -36, 50, -11, 5, -9, 22, -5, 34, -12, -14, 36, -34, 27, 0, 4, 39, -20, 13, -2, 24, -2, 25, -20, -14, 11, 8, -17, -6, -21, -2, 7, 71, -41, 23, 21, 18, -27, -3, 33, 40, -9, -16, 24, -55, 25, -4),
    (-22, 8, -15, -43, 12, 37, 15, -25, -36, 41, 46, 41, -61, -35, 3, -8, -16, -73, 15, 16, 13, 13, -9, 12, -38, 20, -42, 16, 7, -11, -43, -45, -48, 53, 23, 57, -55, 8, 50, -30, -47, 87, 38, 20, 12, -5, -9, -29, 24, -23, -5, 53, 35, -15, -37, 28, -12, 24, -38, -19, 24, -1, 3, -6, -32, 60, -13, 50, -25, -51, 15, -68, -8, -4, -20, -23, -16, -3, -27, -26, 59, 13, -23, -12, 15, -28, 11, 8, 58, -14, -33, -72, 6, 12, 26, -9, 17, 0, 6, 38, -4, 34, -91, -30, -8, -8, 24, -8, -14, -22, -19, -9, 61, 6, 10, 6, 55, -20, -43, -40, 53, 32, 24, 11, -8, 16, -24, -11, -8, 4, 32, 9, -18, 90, 29, -42, 6, -9, 24, -7, -60, -15, -35, -2, 91, 13, 2, 17, 11, 33, -9, -36, 60, 58, 1, 37, 45, 4, -24, -14, -24, -24, 2, -19, -5, 57, -5, -52, 22, 0, -17, 27, 33, -34, 6, -23, 77, 17, -17, 23, -14, 4, 0, -40, -30, -24, -6, 29, 46, -4, -10, 32, -3, -4, -49, 7, 7, 10, 3, -40, -44, 6, -9, -57, 21, -6, 27, -59, 37, 13, 8, 1, 2, 8, 18, -28, 32, -13, -33, -14, -55, 1, 9, -37, 23, 10, -60, 1, -6, 0, 12, 14, -15, -4, 34, -19, 7, -3, -19, -53, 38, 25, -22, 14, 8, -16, -56, 7, 23, -14, -11, 9, -17, -54, -12, -36, -7, -39, -7, 17, 32, -73, 48, 27, 24, -25, -16, -52, -7, -1, -28, -6, -40, 13, 21, 40, 16, -56, -34, 32, 12, 40, -27, -12, 22, -9, -28, -16, -23),
    (-6, 23, -40, 1, -49, 24, 16, 25, 6, -27, -20, -20, 13, 67, -67, 3, -6, 7, -26, -42, -30, -9, -13, 6, -38, 8, -4, -30, -11, 21, 35, -26, 6, 3, -48, 39, -36, 33, -17, 23, 29, -33, -1, -11, -7, 82, -112, -24, -6, -32, -41, -54, -102, -25, -59, -17, 26, 30, 1, 5, 7, -9, 66, 0, -12, -46, -34, 15, 41, -9, -10, -83, 22, 8, 18, -33, 34, -7, -93, -22, -12, 38, -18, -3, -10, -19, -64, -14, 35, 9, -3, 23, -7, 5, -6, 20, -9, -7, -30, 7, -7, -3, 2, 26, -17, -8, -20, -1, -2, 58, -7, 43, -27, -42, -1, -34, -83, 4, -31, 42, -60, -11, -4, 9, 21, -26, 28, -28, -8, 22, -36, 23, -7, -6, -65, 33, 2, -9, -22, -8, 41, 48, -12, -18, -38, -24, 13, -52, -98, -53, 34, 32, -50, 24, -14, 26, 12, 4, 60, -7, -5, 14, -37, -1, 35, 35, -9, 28, 31, 7, -8, -12, 14, 10, -15, -58, -9, 18, 6, -21, -8, -21, -25, 5, 40, -13, -6, 3, -7, -8, 12, 2, -14, 9, 9, 17, -5, 41, -34, 39, -8, -8, 6, -30, -21, 29, 5, 28, -30, 0, -19, -18, -29, 15, 23, 50, -8, -5, 26, -5, 36, 0, 6, 7, -11, 41, 19, -12, 11, 11, -12, 3, -2, 2, 7, -20, 7, 14, 25, 14, -32, -48, -2, 10, -6, 0, 32, 28, -33, -9, 10, -24, 5, 6, -12, 8, -22, 18, 50, -9, 32, 26, 12, 6, 10, -12, 42, 9, -11, -1, 31, -45, 14, 27, -32, -6, 18, 38, 5, 23, 26, -32, 16, 33, 5, 6, 45, 28, -2),
    (-12, 5, 29, -40, 36, -31, -13, -8, -12, -17, 8, -60, 30, 3, 31, -34, 18, -10, 33, -11, -18, 15, 6, 2, -47, -84, 19, -42, -62, -51, 21, 4, -27, 32, 3, -57, -49, 7, 70, -23, -102, 26, 72, 26, -25, 25, 40, 45, 27, -79, 29, -9, -27, 42, 8, 7, -64, -66, -1, -120, 19, -58, 24, -28, -29, 31, -40, -50, -32, -40, -1, -38, -32, -29, 26, 23, -14, 8, -32, -6, 6, -20, 54, -9, 9, 26, -23, 8, 14, -22, 18, -57, -21, -12, 39, 14, -41, 36, -42, -35, -12, 22, 56, -22, -41, 34, -7, 0, -37, 34, 10, -1, 1, 20, 24, -6, -41, 51, 2, -45, 33, 10, -17, -14, -17, -22, 8, -3, -28, -4, 13, -6, 27, -16, 6, -36, -23, 8, 28, 23, -12, -2, 9, -6, 38, -71, 14, 10, 11, 55, -9, -18, -11, -52, 30, -11, -29, -52, 26, -9, 3, -7, -40, -47, 8, 10, 36, -8, -39, 2, 15, 45, 4, 9, 14, 43, -7, -18, 28, -7, -12, 57, 41, 25, -3, -4, -28, -26, 9, -38, 10, -13, -26, -30, 53, -3, -16, 24, -5, 71, 55, -13, 26, 18, -19, 4, -1, 9, 1, 10, -19, -24, 55, 5, 37, 31, -9, 20, 9, 25, 20, 2, -14, 17, -7, 24, 5, -62, -2, -52, -39, 26, 36, 22, -30, -26, 21, 27, 25, -5, 0, 1, 25, -10, -44, 36, 6, -35, 11, -3, 17, -25, -24, -5, 0, -9, 9, 22, -42, -10, 17, -48, -40, -23, 9, 36, 29, 31, 38, -14, -2, 40, -8, 5, -16, -27, 15, -12, 2, -46, -14, 42, 22, -32, 12, -11, -7, 55, -10),
    (32, -15, 48, 10, 32, -57, -51, -30, 34, 40, -7, -24, 28, -43, 37, -9, -42, 31, 14, 7, 67, 37, 23, 3, -28, -1, -7, 43, 14, 8, 15, 20, -5, 11, 73, -16, 52, -75, -49, -46, -17, 15, -65, -19, 4, -79, 100, -17, -67, 38, -17, 39, 85, -18, 37, 4, 46, -53, -16, 15, -70, -10, -21, 18, -7, 57, 51, -28, -5, -12, -9, -8, 13, -9, -6, 8, 7, -38, 0, -19, -59, 43, -1, 29, 2, -59, 36, 47, 10, -5, -1, 19, -16, -7, -62, 1, -1, 23, 17, 8, 13, -28, -27, -16, 39, -27, -45, -24, 42, -41, 31, -43, -42, 42, 22, -38, 47, 17, 26, 39, 14, 20, -34, -24, 16, -27, -17, 11, -8, 35, 30, -23, 60, -40, -24, -2, 12, 25, -75, -4, 20, -51, 39, -6, -39, 34, 5, 20, 56, 21, 11, 56, 20, -14, 18, -2, -32, -62, -24, 12, 2, 8, 12, 6, 27, -10, 12, -4, 3, 19, -24, -19, -35, -37, 18, -32, -8, 24, 5, 40, 20, 33, 21, 26, -43, -16, -21, -8, -67, 15, -25, 3, 25, 24, 0, 8, -2, -16, 16, 22, 18, 31, -15, 28, -9, -15, 25, 8, -26, -3, -8, 9, -7, -3, 31, 28, -10, 24, -8, -20, 23, 24, -8, -9, 13, 39, 18, 8, -18, 13, -2, 11, 8, 29, -7, 26, 45, -9, -11, 9, -18, 9, 13, -8, -19, 13, 9, -3, -14, 46, -9, 0, 29, 12, 16, -11, 27, -19, -10, -21, -10, 14, 6, 16, 24, -18, 6, 31, 26, 11, 15, -13, -8, 24, 48, 7, -10, 31, 15, -11, -30, 42, -16, 17, -15, -10, -12, 25, -13),
    (-2, 7, 24, -6, 10, -30, 19, -9, 41, 9, -10, 21, 32, -23, 10, -32, -13, -49, 24, -29, -39, -9, 1, 13, -94, -7, 3, -2, 40, 17, 11, -9, 37, -16, 8, 37, 51, -64, -8, -37, 10, -21, 2, -44, 40, -22, -11, -41, -98, 48, 23, -8, 4, 31, 1, -13, -23, 2, 7, -12, -34, 2, -21, 19, -46, -35, 6, 4, 31, -36, -9, -52, 10, -57, -21, 0, 16, -101, 63, -9, -82, -6, -3, 7, 59, 0, 30, -10, -3, -9, 8, 7, -47, -19, -45, -26, -48, 27, -4, -51, 11, 27, 18, 1, -26, 17, 17, 16, 74, -2, -58, -31, 23, 3, 62, -39, -63, -27, -1, -19, -13, -22, -21, 4, 59, 17, -7, 36, 21, -49, -9, 8, 33, -43, 21, -28, 38, -25, -28, -31, 49, -43, -4, -40, -74, 12, 7, 29, 43, 33, 52, 35, -24, -13, -49, 39, -18, 40, 24, 7, -66, 26, 39, 8, -20, -11, -37, 40, 9, 20, -32, 28, -27, -73, 28, 5, -38, -44, 6, -7, 26, 4, 25, 27, -5, 3, -22, 36, -42, 20, -48, -33, -21, -15, 3, -19, 67, -48, -8, -7, 22, -21, -25, -18, 71, 24, -69, -2, -3, 14, 25, -36, -45, 11, 2, 15, -11, 21, -19, -9, 11, -2, 12, 13, -8, -29, 22, 3, 26, 11, -18, -15, -2, -11, -24, -7, -2, -27, -17, 14, -36, 5, 20, 57, 31, 40, 38, 20, -31, -5, -47, 43, -22, -3, 4, -13, -56, -10, 66, -22, 17, 3, 31, 22, 31, 32, -3, 49, -8, 4, -18, -5, -34, 35, 11, 19, 67, 0, 33, 31, -44, 15, 26, -19, 34, 28, -15, 1, -9),
    (-24, 12, 0, -19, 38, -26, 8, -16, -3, 31, 19, 41, 3, -23, 55, 25, -37, -69, 37, 42, 6, 35, 39, 46, -41, -17, -9, -32, -23, 40, 3, -2, -32, 61, -8, -58, 41, -34, -11, -5, -5, 30, -14, -1, -12, -24, 23, -34, -20, -58, 46, 1, 22, 100, 53, 11, -41, -75, 38, -46, -22, 25, 15, 48, -19, -20, 54, -41, -40, -9, -31, 32, 15, 30, -9, 5, -23, -16, 42, -19, -41, -20, 8, -13, 22, 46, 70, 13, -38, -17, 24, -46, -33, 20, -36, 10, -4, 28, -52, -8, -70, -51, -29, 7, 21, 14, -2, 33, 7, 52, 16, 7, 12, 15, -8, 5, -48, -71, -19, 21, 9, -62, -27, -33, 7, 25, -17, -13, -20, -20, -4, -17, 6, -41, -34, 39, -2, 36, 28, 31, 13, 45, -11, -9, -8, -25, -55, -19, -78, -75, 4, -43, 1, -9, 32, -37, 26, 17, 12, -30, -57, -6, -10, -9, 11, -56, -15, 53, -17, 29, 33, -10, 33, 9, -15, 9, 45, -38, 1, 13, -47, -64, -50, 13, -8, 28, 31, 6, -4, 44, -19, -20, -64, 6, 12, -42, 11, -18, -3, 41, -20, 31, 26, 2, -23, -33, 9, 22, 18, -12, -45, -2, -5, -47, 19, -62, 6, 27, 70, 24, -17, -15, 14, 66, 7, 3, -13, 23, 27, 22, 27, -17, -4, -23, 25, 7, 26, -1, 14, -7, -47, -2, -25, 70, -20, 9, -31, 35, -2, 69, -46, 40, 0, -11, 30, -55, -4, -17, 29, 34, 30, 27, 29, -44, -7, -30, 0, -7, 3, 7, 53, -28, -33, 33, -38, 15, 37, -12, 5, 22, 11, 10, -40, 26, 15, 20, 69, -66, 12)
  );
  ----------------
  CONSTANT Flatten_1_Columns : NATURAL := 2;
  CONSTANT Flatten_1_Rows    : NATURAL := 2;
  CONSTANT Flatten_1_Values  : NATURAL := 32;
  ----------------
  CONSTANT NN_Layer_1_Activation : Activation_T := relu;
  CONSTANT NN_Layer_1_Inputs     : NATURAL := 128;
  CONSTANT NN_Layer_1_Outputs    : NATURAL := 10;
  CONSTANT NN_Layer_1_Out_Offset : INTEGER := 6;
  CONSTANT NN_Layer_1_Offset     : INTEGER := 0;
  CONSTANT NN_Layer_1 : CNN_Weights_T(0 to NN_Layer_1_Outputs-1, 0 to NN_Layer_1_Inputs) :=
  (
    (-1, -79, 4, -74, -107, -20, -64, -40, -44, 4, 33, 110, -47, -53, 32, 35, 41, 10, -48, 64, -33, 7, 56, -21, -6, 52, -4, 105, -69, 32, 42, 33, 18, -31, -47, -41, -52, -18, -57, -25, -44, -24, -20, 12, -27, -4, 36, 20, -17, -4, -4, 12, -8, -26, 23, 44, 1, 55, -18, 4, 19, 32, 7, -47, 23, -56, -53, 22, -49, -11, -14, -35, 6, 17, 14, 25, -4, -55, 3, 2, -20, -13, -43, -3, 33, -11, 26, -7, -5, 19, -31, -20, -40, 3, -19, -17, 12, 22, -10, -13, -7, 2, -12, -26, 15, 5, 13, 9, -13, 3, -1, -5, -16, 6, 4, -7, -21, -17, -14, -5, -5, 16, -30, 13, -9, 13, 21, -19, 17),
    (32, -10, -92, -39, -55, 32, 0, -32, 32, 27, 55, -20, 4, 69, 11, 1, 58, 39, -12, -14, -11, -39, -20, -21, 28, -48, -38, 24, -4, -44, 16, -22, 14, -38, -62, -22, -52, 13, -18, -15, -4, 9, 27, 16, 5, 53, 27, -5, -4, -4, -12, -2, 9, -9, -1, -15, 35, 12, 11, 11, 45, -36, -44, -26, 14, 26, 1, -21, -28, 21, 7, -17, 26, -13, 24, -15, 12, -5, -40, -12, 18, -9, 14, 19, 8, -16, 10, -9, 43, 5, -10, 11, 8, 31, 19, -2, -1, 26, -4, -19, 12, 41, -13, -31, 16, 10, 33, -9, -15, 39, -17, -16, 2, 22, -9, -14, 15, 7, -33, 4, 5, 13, 9, 17, -46, 7, 11, 8, 19),
    (-26, -47, -11, 38, -19, -28, 40, 12, 4, 22, -61, 2, 32, 28, 62, -48, 18, -50, -2, 4, 23, -9, 12, 7, -43, -62, -7, 78, 4, -48, -32, -35, 4, -20, -16, 35, -12, -16, -5, -2, -23, 32, -9, 13, 6, -32, -17, -22, -20, -53, -14, 20, 14, -40, -2, 0, -38, -30, -34, 21, -23, -44, 6, 18, -15, -27, -21, 43, 7, -10, 29, 11, 30, 28, -9, -19, -4, 40, 12, 0, 22, -36, -6, -1, -21, 2, -11, 4, 21, 0, -11, -10, 22, -3, 5, 35, -2, -47, -7, 6, -18, 1, -8, 11, -6, 3, 1, 1, 3, 4, 6, 5, 13, -1, 12, 19, 21, -5, -7, -4, 8, -6, -7, 23, 8, -21, 15, 22, -4),
    (-56, 56, 11, 35, 63, 42, -43, 9, -28, -39, 47, -78, -76, -4, -3, -63, 0, -29, 44, -16, -4, 8, 63, -50, 42, 27, 32, -2, -58, 19, 21, -16, -15, 8, -35, 4, 8, 9, -16, -35, -24, -7, 23, -23, -5, 3, 8, 16, 12, 1, 12, -13, 15, -7, 5, -12, 14, 46, -12, 5, -9, 19, -3, -16, -4, 41, 8, 29, 28, 26, -5, 34, -64, -49, 0, -12, -32, -66, -2, 17, 8, 28, 15, -44, -2, -18, 17, -38, 4, 6, 2, 14, -23, 9, 5, -57, 19, -3, 5, 12, 2, 27, 2, -16, 11, -5, 1, 0, -49, -1, 5, -22, 1, -16, 25, -43, -19, -32, 18, -37, 9, 14, -3, 6, -24, 41, 1, -16, -18),
    (30, -17, 22, 40, -26, 27, 16, 37, -14, -44, -53, -42, 36, -2, 7, 1, -108, -64, -6, -13, -14, 36, -39, 47, -65, 11, -29, -41, 2, 36, 21, 63, -21, 10, 57, 1, 11, 28, 20, 17, 46, -51, -23, -13, 30, -20, -24, 2, -13, -47, -15, -16, -10, 2, 15, 21, 22, -52, -27, -37, -43, 57, 26, 22, 5, -21, -5, 59, -12, 18, 14, 10, 16, 8, -24, -8, 5, 25, 7, 14, 31, -64, -16, 10, -3, -18, -40, -9, 14, -6, -25, -18, 39, -28, -1, 19, 5, -27, 3, -2, -14, 12, 1, 11, 6, 15, 4, 8, 14, 24, 33, 11, 17, -17, -9, 7, -9, 11, 14, 12, -23, -11, 4, 14, 1, -15, 1, 19, 13),
    (-21, -49, 1, -39, 60, -6, -108, -51, -93, -54, -22, -28, 29, 40, -48, -44, -33, 32, -25, -25, 28, -8, -41, 11, 25, 20, -43, -44, -58, 76, 55, -8, 7, -56, 22, -18, 20, -15, -36, -18, 5, -46, 18, -10, 29, 11, -35, 4, -12, -26, 14, -10, -9, -21, 19, 30, 14, -13, 2, -36, -1, 34, 18, -7, -34, -21, 31, -15, 73, -40, 1, -36, -34, -23, -43, 12, 36, -10, 9, -15, -25, -14, 5, 18, -6, -4, -53, 3, 5, -20, 11, -38, -1, 37, 42, 9, -10, 29, 6, 14, 34, -4, -9, -25, -14, 12, 7, 5, 16, -12, 3, 16, 2, 29, -23, 36, 0, -3, -26, -15, 7, 3, 27, -15, -24, 15, 22, 1, -34),
    (20, 25, -19, 23, -36, -9, 34, 43, 43, 4, 6, -24, -62, -43, 18, 46, 51, 67, -27, 48, -74, -51, 33, -68, -60, 3, 36, 8, -21, -83, -95, 22, -13, 3, 26, -24, -28, -23, 4, 44, -7, 6, 9, 8, -28, -13, -14, -3, 49, 35, 9, 18, -11, -1, 18, -5, -20, -35, 11, -12, 16, -47, -1, -32, 19, 28, -18, 26, -49, 20, 4, 23, 37, -5, 8, -22, -13, -50, -19, -5, 2, 3, -15, -58, 14, -2, 37, -2, -29, 26, -8, -3, -43, -13, -16, -22, 34, 7, -3, -26, -15, 14, -32, 2, 4, -13, -33, -4, -14, -26, -26, -17, -23, 30, 19, -10, -24, -38, 33, -39, 3, -10, -27, -21, -11, 12, -4, -23, -34),
    (-15, 23, 28, -12, -13, -19, -21, -20, -28, 50, 3, 19, 32, -6, -10, -20, 10, 27, 44, -32, -25, 43, -39, 24, -50, -9, 20, 28, 4, 11, 17, -32, 7, 31, -3, 13, -4, 24, -22, -16, 10, 26, 0, 7, -1, 3, -14, 6, -4, -20, 15, -4, 14, -4, 6, 9, -26, 1, -1, 10, -12, 2, 10, 22, -11, -6, 4, 4, 9, -15, -4, -33, -1, 30, -42, -12, 39, 13, -21, -14, -11, -4, 34, 41, 2, 18, -5, 30, 12, -35, -9, -28, -20, 3, 17, 28, 12, -3, 16, -6, -5, 6, 0, 7, -37, -8, 21, 17, -10, -19, 9, -8, 13, 9, 22, 12, -4, 9, -24, 16, -17, -36, -7, 6, 6, -13, 13, 15, 24),
    (-5, 35, 22, 28, 59, -4, 41, 2, -11, 24, -27, -57, -80, -38, -46, -48, -33, 0, 59, 2, 0, 17, 25, -6, -4, -63, 52, -30, 18, -3, -44, 27, 5, 10, 10, 10, 15, -9, 3, 21, 10, 27, -30, 9, -16, -29, 9, 11, -25, 44, 1, -15, -19, -34, 2, -19, -9, -62, 35, 3, 4, -24, -11, 10, 23, 38, -3, 20, 17, 9, -1, 40, -1, 5, 8, -13, -36, -38, -5, 34, 3, 13, -9, -56, -3, -1, 31, -25, 0, 26, 29, 30, -3, -26, -35, -26, -6, -17, 20, 18, -13, 7, 4, -6, 10, 11, 18, 3, -20, -4, -32, -4, -14, 7, -10, -12, -2, 5, -8, 1, -5, -15, -11, 3, 8, -18, -9, -37, 19),
    (54, 7, 5, -94, 14, -41, 40, -43, -20, -14, 2, -11, 4, 32, -70, 33, -24, 35, -86, 79, 37, 36, -97, -53, 36, -10, 4, -30, -7, -10, 14, -4, 4, -18, 45, 7, 11, -33, 32, 29, -17, -41, 42, 29, 18, -19, -26, 31, -25, 2, 23, 27, -27, 18, 11, -46, -19, 36, 17, -24, -18, -29, 37, -8, -34, 3, 21, 1, 44, -54, 12, -37, 18, -25, -36, 26, 27, 1, -11, -14, -24, -13, 4, 1, 27, 11, -3, 22, 10, -12, -42, -21, 21, 10, -18, 31, -19, 11, 0, -3, 29, -12, -1, -24, -8, -8, -15, -18, -25, 18, 22, 30, 9, 8, -15, 10, 12, 26, -20, -2, 22, 10, -3, -18, 22, 3, 3, 7, -1)
  );
  ----------------
END PACKAGE CNN_Data_Package;
