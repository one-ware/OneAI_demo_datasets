library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.numeric_std.all;
use work.CNN_Config_Package.all;

PACKAGE CNN_Data_Package is
  CONSTANT Layer_1_Columns    : NATURAL := 128;
  CONSTANT Layer_1_Rows       : NATURAL := 128;
  CONSTANT Layer_1_Strides    : NATURAL := 1;
  CONSTANT Layer_1_Activation : Activation_T := relu;
  CONSTANT Layer_1_Padding    : Padding_T := same;
  CONSTANT Layer_1_Values     : NATURAL := 1;
  CONSTANT Layer_1_Filter_X   : NATURAL := 3;
  CONSTANT Layer_1_Filter_Y   : NATURAL := 3;
  CONSTANT Layer_1_Filters    : NATURAL := 12;
  CONSTANT Layer_1_Inputs     : NATURAL := 10;
  CONSTANT Layer_1_Out_Offset : INTEGER := 3;
  CONSTANT Layer_1_Offset     : INTEGER := 1;
  CONSTANT Layer_1 : CNN_Weights_T(0 to Layer_1_Filters-1, 0 to Layer_1_Inputs-1) :=
  (
    (-20, -11, 17, -1, 53, 38, -17, 27, 17, 0),
    (4, -15, -48, 0, -29, -6, 24, 15, 58, 0),
    (-18, 20, 10, 41, 33, 49, 25, 38, 12, -2),
    (7, 68, 22, 17, 14, 12, -22, 3, -39, 0),
    (-1, 41, 31, 31, -50, -3, 13, 22, 21, 3),
    (22, -5, 11, 46, 17, 37, 22, -30, -31, 1),
    (-29, -23, -26, -14, 11, -9, 34, 39, 13, 0),
    (33, 20, 38, -8, -3, -14, -23, -26, -36, -1),
    (42, 0, -12, 3, 35, -41, 14, -16, -38, -1),
    (26, -15, -7, -33, -25, -22, -7, -23, 44, 3),
    (46, -10, 31, -7, -26, -7, 1, 7, 40, -5),
    (54, -34, -47, 26, 10, -44, -19, -62, -45, -3)
  );
  ----------------
  CONSTANT Pooling_1_Columns      : NATURAL := 128;
  CONSTANT Pooling_1_Rows         : NATURAL := 128;
  CONSTANT Pooling_1_Values       : NATURAL := 12;
  CONSTANT Pooling_1_Filter_X     : NATURAL := 2;
  CONSTANT Pooling_1_Filter_Y     : NATURAL := 2;
  CONSTANT Pooling_1_Strides      : NATURAL := 2;
  CONSTANT Pooling_1_Padding      : Padding_T := valid;
  ----------------
  CONSTANT Layer_2_Columns    : NATURAL := 64;
  CONSTANT Layer_2_Rows       : NATURAL := 64;
  CONSTANT Layer_2_Strides    : NATURAL := 2;
  CONSTANT Layer_2_Activation : Activation_T := relu;
  CONSTANT Layer_2_Padding    : Padding_T := same;
  CONSTANT Layer_2_Values     : NATURAL := 12;
  CONSTANT Layer_2_Filter_X   : NATURAL := 3;
  CONSTANT Layer_2_Filter_Y   : NATURAL := 3;
  CONSTANT Layer_2_Filters    : NATURAL := 16;
  CONSTANT Layer_2_Inputs     : NATURAL := 109;
  CONSTANT Layer_2_Out_Offset : INTEGER := 3;
  CONSTANT Layer_2_Offset     : INTEGER := 0;
  CONSTANT Layer_2 : CNN_Weights_T(0 to Layer_2_Filters-1, 0 to Layer_2_Inputs-1) :=
  (
    (0, -6, 9, 18, 1, 26, -45, -68, -37, -39, -16, -43, 17, -28, -18, -4, -4, -4, -23, -19, -40, -53, 21, -40, 7, -49, 8, -10, -15, 17, -48, 0, -32, -44, -15, -10, 23, -6, -19, 13, -5, -6, -69, 9, -21, -26, -19, -22, -32, -50, 24, 20, 14, -13, -73, 18, -18, -23, 4, -5, -24, -31, -10, 15, -9, 28, -66, 15, 3, -2, 5, -1, -2, 11, 8, 6, 17, 38, 7, 25, 9, 17, -25, 0, -19, 25, -7, 26, -6, 26, 17, 8, 37, 17, -7, 22, 6, 4, 7, 22, -19, 7, -14, 8, 32, 28, 2, 18, -4),
    (-9, -48, -22, 27, 13, 42, -38, 33, 39, 6, 22, -19, -17, 14, -24, 23, -14, -19, -6, -1, 13, 22, -20, -51, 7, 0, -26, -9, -22, 2, 27, 39, -15, 13, -15, -26, -38, 10, 2, 11, -4, -26, 14, 32, 6, 23, -28, 22, -21, -5, -8, -25, 6, -20, 24, -23, -26, 16, -16, -14, 3, 27, 16, -14, -28, 0, 34, -9, -79, 16, -11, -56, -12, 16, -8, -23, -5, -15, 16, -39, -30, -12, -18, 46, 5, 0, 30, 6, 16, -8, 20, -9, 3, 12, 10, -39, 20, 24, 40, -6, 30, -7, 30, 8, -22, -2, 20, -57, -2),
    (-5, 22, -10, -22, -4, 18, 5, -28, 1, 13, -21, -30, -4, -20, 9, -10, -15, -10, -9, 11, -16, 0, -53, -55, -12, -34, 19, 12, -17, -7, -1, -3, -17, -17, 13, -10, 8, 10, -1, -9, -9, 29, 25, -58, 27, 2, 14, 3, -18, -12, -4, -32, 14, 7, 12, -40, 29, 3, -2, 14, 1, -26, 8, 16, -5, -21, -22, -11, -14, -26, 6, -10, -14, -2, 15, -26, 37, 28, 28, -21, 10, 0, 38, 0, -7, 12, 9, -34, -21, 7, -29, -28, 23, -11, -24, -17, -29, -12, 8, -11, 1, 3, 1, 15, -13, -20, -9, -26, 1),
    (34, -1, -15, 10, -10, 13, -16, 9, -27, 12, 5, 59, 9, -19, -3, 13, -7, -3, 21, 3, 15, 23, 26, -1, 18, -8, 28, 12, 14, 12, 13, 6, -9, 9, 27, -4, -6, -28, -2, 29, -17, -4, -33, 45, 9, 12, -6, 14, -7, -23, 20, 11, -11, 1, -21, 49, -23, 16, 10, 1, -21, -2, -19, 27, 16, 37, 17, 26, -2, 25, -8, -19, -3, 20, -1, -12, -1, -36, 42, 30, -17, 11, -29, -1, -33, 24, 0, -45, -2, -43, 27, 18, -13, 12, -13, -46, -18, 26, -22, -22, -40, -27, 47, -32, -48, 3, 4, -41, -2),
    (36, -18, 31, 7, -37, -13, -16, 7, 13, 20, -19, 67, 32, -12, 12, 9, -35, -11, -22, -17, 11, 22, 7, 49, 5, -12, 27, -3, -7, -17, -1, -1, -6, 31, 3, 25, 28, -10, 21, -11, -13, -14, 31, 10, 45, 35, -1, 60, 26, -12, 4, 34, -25, -3, 16, 0, 39, 44, -3, 43, 26, -6, 26, 2, -27, 3, 5, 10, 30, 16, 14, -11, 6, -10, 2, -6, -1, 18, 12, -25, -9, 31, -11, 16, 16, -7, 5, 32, -13, -5, 24, -8, 25, 20, 4, 6, 36, 16, -8, 8, -16, -3, -13, -3, 9, 3, 13, 6, -3),
    (-41, -18, 7, -39, -2, -3, -40, -40, -6, 8, -17, 29, -12, 8, 2, -22, -17, -16, -1, -69, -13, 21, -21, -31, 1, -9, 1, 7, 18, 2, -4, -19, 19, 35, 5, 54, -9, -18, 5, -51, -7, 2, -6, -33, -19, 26, -22, 2, 16, 15, -12, 15, 9, -28, -27, -36, 17, 11, 7, -14, 36, -10, -16, 15, 35, 8, 11, -27, 17, 56, 27, 75, -15, 3, -27, -29, -25, -3, -19, -18, -26, -7, -18, -5, -6, -2, -11, 27, -13, 4, 9, -46, 12, 26, 8, -44, 8, 26, 31, -16, 15, 15, 26, -15, 28, 6, 35, 37, -1),
    (-11, -2, -8, -18, -21, -28, 7, -2, -20, -10, -25, -40, -12, -20, 18, -9, 23, -8, -8, -37, -16, 0, -4, -11, -24, 11, -9, 15, -13, -14, 0, -42, 8, 13, -8, -9, 0, 5, -2, -5, 14, -13, -19, -26, -22, 28, -13, 4, -6, -33, -9, -17, 24, 8, -9, -23, -21, 27, 16, -30, -17, -10, 11, -24, -8, 35, -21, 1, -16, 1, -8, 12, 21, -23, -43, 7, -11, -36, -21, 5, -12, -12, -30, -31, 2, 3, -30, -18, 14, -41, -32, -13, -7, 4, 1, 16, -25, 36, 7, -10, 4, -29, -4, 18, -46, -3, 4, 0, 8),
    (31, 11, -5, 16, 28, 29, -9, 28, 21, 44, 19, 51, 4, -14, -21, -2, 7, -9, 9, 17, 53, 7, -11, 51, -8, 7, 11, 7, -39, -1, -19, -7, 22, -20, -4, 8, 9, -6, 3, 20, 7, 34, 13, 21, 12, 33, -2, 76, -10, -14, -4, 19, -23, 12, -37, 22, 1, 13, 1, 38, 7, -24, 2, 14, -21, -23, -40, -21, -21, 41, -32, 3, -7, 5, -7, -1, 3, 39, 1, 23, -1, 14, 11, 45, -40, -14, -15, -1, -11, 16, -24, 16, -18, 11, 9, 35, -18, 25, -7, -43, -3, -41, 2, -11, -30, -17, -10, -15, -1),
    (-20, 0, 22, -3, -30, -30, 15, -29, -22, -28, 1, -49, 16, 6, 10, 22, -18, 3, 16, -6, -32, 7, -9, 9, 9, -5, 0, 2, -27, -15, -16, -29, -27, -17, 2, 2, 16, -12, -12, -11, 7, -15, -7, -28, -8, -28, 14, -6, -25, -6, 14, -12, 15, 10, 8, 4, 0, -29, -30, -37, 5, 11, -20, -9, -32, -8, 3, -10, 17, 13, -28, -25, -15, -14, -27, 28, -21, -40, -11, 12, -9, -17, -23, -13, 34, -11, 9, 28, 5, -13, 9, 16, -2, -21, -25, -41, -15, -26, -13, -2, -21, -27, -28, -7, -15, 21, -13, 24, -1),
    (-4, -20, 43, 26, 23, 10, -10, -11, -8, 20, 9, 13, -17, 9, 32, 29, 14, -14, -12, -16, 1, -7, 18, -5, 7, -11, 4, 11, 45, -19, -18, 11, -25, 13, 18, -18, 20, 0, 34, 2, 20, 3, 2, 8, 6, -29, -3, -3, 10, 2, 0, 3, 9, 10, 0, 2, -9, -17, -9, -47, 4, 5, 17, 2, 30, -6, -19, 15, -45, 9, 3, -26, 19, 22, -26, -8, -15, 24, -1, 11, -14, -14, -20, -18, -13, 18, -9, 12, -9, 18, -6, 14, -12, -24, -37, -4, -8, -3, 27, -6, 10, 18, 27, 15, -10, 27, -14, -7, 1),
    (-6, -12, -9, -9, 2, -14, 25, 34, -7, -9, 11, 4, -21, -33, -19, 16, 11, -16, -8, 30, 2, -16, -14, 9, 0, -37, 1, 37, 16, 26, -30, 49, 32, -1, 5, -14, -5, 35, 27, -30, -18, 3, 42, 2, 22, -33, -15, -18, -17, 39, 14, -31, -31, -24, 21, 14, -29, -11, -22, -15, 8, -8, -18, 2, -19, -40, 9, 3, -23, 30, -9, -18, 31, 36, 12, 20, 12, 21, -14, 5, 8, -16, 18, 2, 8, 22, 13, 4, 26, 6, 19, -9, -7, 16, -6, -24, -7, 24, 1, -33, 18, -4, 32, -19, -2, -2, -7, -14, -1),
    (-21, -4, -6, 30, 21, -7, -11, -5, 39, 7, 20, 28, -6, -27, 16, 32, 36, 7, -11, -24, 21, 12, 38, 24, 4, -10, 43, 8, 41, -14, -12, 9, -4, 8, 30, -26, -22, -10, 18, 19, -7, 8, -11, -7, 26, -1, -17, 15, 14, -3, 3, -1, 14, 11, -8, 5, -8, 9, -22, 23, -12, 4, -18, 17, 6, -11, -35, -7, 4, -2, -2, -32, -4, 2, 18, 28, 7, -24, 6, 4, -8, -20, -10, -10, 13, -9, -31, 38, 17, -16, 17, -24, 30, -1, -4, 19, 15, -12, 21, 14, -5, 12, -12, -5, -6, 5, -10, 31, -2),
    (16, 7, 6, -23, -34, 21, 48, -3, 33, 9, -8, -23, 37, 22, -5, 4, -28, -24, 32, 12, 28, 29, -23, -11, -2, 25, -12, -6, -30, 7, 10, 23, 20, 1, -29, -9, 4, 2, -7, 25, 8, 24, 47, 18, -2, 27, -30, -18, 36, 18, 26, -20, -24, -2, 34, 13, 19, 48, -27, -12, 37, 20, 27, -4, -27, 14, 16, 3, -14, 26, -8, -17, -14, 1, -5, 4, 15, 23, 34, 19, 25, -9, -1, -9, 15, 22, 17, -21, -25, 5, 20, 20, 5, 20, -21, -8, 37, 37, 14, 4, -2, -15, 5, 3, -20, 27, -7, -34, -1),
    (-5, 2, 25, 35, 2, 7, -1, -7, 10, 5, 13, 22, 6, -3, 19, 33, 11, 21, -48, -11, -4, 31, 24, 45, 1, -22, -11, 21, 13, -22, -60, 29, 41, 3, -11, 13, -11, -42, 29, -22, 7, -4, -29, 13, -15, -10, -30, 10, -29, -20, 21, 15, -15, 26, -21, -20, 1, 17, -8, -31, 1, 20, -18, -23, -21, -44, 18, 7, 11, 3, -27, -13, -19, -8, -21, -21, -28, -17, -11, -9, 8, -12, 3, 9, 19, 12, -12, -37, -45, -25, 15, -35, -10, 11, 3, -3, 21, 10, 11, -16, -2, -11, -14, -52, -92, 0, 29, -75, -3),
    (-13, -45, 13, 14, 10, 4, 1, -14, -36, -36, -16, 4, -55, -45, -17, 46, -12, -13, -57, -4, 25, -15, 30, 11, 12, 21, -9, -1, -10, -17, -7, 0, -8, 13, -16, 20, -28, -16, -33, -26, -32, -3, 14, -7, -36, -28, -21, 5, 8, 15, -2, -15, 3, -7, 17, -25, -20, -15, 20, -60, -7, 24, -18, -29, -1, 36, 12, -11, -66, -6, 16, -24, -12, -11, -31, -23, -33, 8, -29, -4, -5, 10, 1, -36, 5, -1, -8, -9, -12, 26, -26, -13, -6, -40, 6, -15, 18, 12, -6, -7, -14, 23, 23, 13, -50, -29, 2, -36, 0),
    (11, 21, -12, 3, 5, 39, -14, 3, 3, -17, 6, 18, -7, 18, 21, -3, 25, -17, -13, -32, 21, -14, 1, -26, -1, 24, 4, -21, -26, -7, -16, -18, -17, -21, -8, 31, -13, 22, 29, 16, 26, 28, -5, -31, -23, -11, 23, 6, 18, 14, 3, -16, 43, -6, -8, -31, 1, -21, 15, -16, -9, 10, 7, 5, 5, -9, -13, -33, 5, -9, 3, -9, 1, 23, 34, -13, 21, 23, 12, -41, -6, -31, 30, 9, 17, 28, -7, -23, 17, -20, -4, -23, -25, -42, 5, 2, 22, 24, -6, -8, 39, -15, -28, -35, -29, -21, 31, -25, 1)
  );
  ----------------
  CONSTANT Layer_3_Columns    : NATURAL := 32;
  CONSTANT Layer_3_Rows       : NATURAL := 32;
  CONSTANT Layer_3_Strides    : NATURAL := 2;
  CONSTANT Layer_3_Activation : Activation_T := relu;
  CONSTANT Layer_3_Padding    : Padding_T := same;
  CONSTANT Layer_3_Values     : NATURAL := 16;
  CONSTANT Layer_3_Filter_X   : NATURAL := 3;
  CONSTANT Layer_3_Filter_Y   : NATURAL := 3;
  CONSTANT Layer_3_Filters    : NATURAL := 24;
  CONSTANT Layer_3_Inputs     : NATURAL := 145;
  CONSTANT Layer_3_Out_Offset : INTEGER := 3;
  CONSTANT Layer_3_Offset     : INTEGER := 0;
  CONSTANT Layer_3 : CNN_Weights_T(0 to Layer_3_Filters-1, 0 to Layer_3_Inputs-1) :=
  (
    (1, 28, -32, -19, -10, 10, -5, 2, 29, -14, -31, -21, -10, -2, 18, -14, 22, 59, -61, -12, 14, 18, 10, 19, 2, -9, -37, 3, -3, 10, 30, 15, 7, 27, -35, -5, 2, 20, 12, 7, 20, 6, -9, 19, 7, -2, -14, 17, 30, 46, -36, 11, 8, 21, -3, 25, -19, 22, -36, 13, -14, 9, 2, 4, 39, 70, -33, -2, -4, 41, -28, 41, 1, -1, -54, -10, -27, 28, 7, 13, 27, 40, -25, -14, 1, 7, 35, 23, -1, -3, -28, 2, -14, 33, -5, -2, 25, 24, -25, -3, -18, 4, -22, 26, -1, 24, -21, 7, -7, 17, 20, -1, 20, 43, -14, -9, -5, 17, -17, 24, 18, 7, -30, 13, -20, 19, 1, 1, 35, 30, -21, 2, 8, 6, 22, 13, -3, -23, -17, -10, -9, 12, 21, -21, -2),
    (20, -4, 12, 32, -21, -15, -1, -55, 25, -13, 20, -25, 3, 21, 18, -5, 35, -21, 37, 32, -27, -28, -9, -46, 0, 0, 48, -19, 6, 0, 37, -10, 3, 2, 6, 28, -6, -14, 22, -49, -17, 4, 22, -16, 8, 7, 27, -5, 12, -5, -15, 15, -17, -29, 9, -15, 22, -5, 25, -28, 14, 29, 3, -1, -1, -9, 2, 31, 2, -33, -30, -49, -10, 14, 43, -25, 16, 21, 3, 13, 13, -1, -2, 31, -13, 7, 3, -29, 10, 4, 24, 2, 25, 17, 13, 17, -9, -3, -41, 4, 16, -1, -10, -7, -33, -11, 17, 13, 5, 6, -14, -28, 22, 8, -4, 12, 16, -7, 1, -24, 2, -18, 22, -14, 9, 39, 4, 15, 24, 7, 8, 4, -12, -25, 0, -11, -29, 25, 18, 4, -1, 23, 2, 15, 2),
    (11, 7, -51, 22, -9, -9, -58, 22, -43, 18, 12, 15, -14, 11, -21, 12, 18, -5, -11, 39, -8, -12, -14, -2, -2, -6, 22, 3, 13, 26, -31, 0, -4, 8, -5, 35, 20, -13, -36, -14, -23, 27, 7, 1, 5, 7, -2, -8, 19, 0, -20, 22, 4, -17, -16, -2, 13, -17, 23, 18, -1, 23, -16, -11, 31, 7, -10, 51, 17, -30, -43, -17, -9, 1, 30, 2, 10, 32, -18, -25, 13, -4, -10, 37, 11, -19, -41, -18, 7, 10, 16, -4, 6, 28, 12, -18, -1, -21, 13, 1, -8, -2, -19, -3, -24, -17, 28, 11, 11, 19, -10, -29, 15, 19, -3, 28, 21, -20, -19, -3, 33, 17, 16, -19, 17, 14, 16, 0, 19, 29, -3, 7, -8, -24, 1, 20, 16, -6, -5, 6, 8, 34, 0, -29, -1),
    (12, -6, 4, 19, 11, -23, -26, 3, -31, -2, 9, -21, 9, 9, 4, -27, 0, -17, -28, -12, 37, -4, -6, 2, 9, 3, 3, -13, 31, -23, -18, -22, -8, -2, -13, -10, 17, 4, -19, 2, -8, -8, -2, 2, -5, -1, -1, -21, -1, 2, 2, 8, 13, -4, 4, 10, -3, 7, 8, -21, 36, 17, -9, 1, 2, 19, -30, -3, 31, 8, 10, 14, 12, -16, -12, -4, 48, 10, 1, -7, -1, 17, -1, -5, 32, 10, 8, -1, -32, 3, -16, -9, 24, 1, -14, -17, -3, 1, 32, -1, 4, -15, 7, -7, -6, 7, 21, -3, 25, -16, 20, -6, 2, 18, -19, 2, 31, -4, -11, -1, 7, 10, 14, -6, 6, -19, -24, 1, 11, 21, 1, -3, 22, 29, -17, -8, -34, 7, -3, -22, 10, 4, 17, 9, -2),
    (-1, -32, 46, -37, 18, 19, -15, 5, -14, -3, -17, 26, -18, -29, -23, 3, -8, -8, 27, -19, 22, -23, -30, 6, -4, 9, 7, -1, 20, -26, 14, 13, 4, 35, 7, -14, -4, -1, 51, -9, -8, -3, -8, 18, 25, 13, 38, 34, -13, -37, 20, 7, -26, 7, 10, -8, 18, 15, -27, -20, -24, -1, -34, 8, 0, -29, -8, 15, 5, -32, -14, -32, 23, -8, -7, -18, 4, 1, -17, -2, 35, 29, 13, 24, 5, -33, 24, -18, 13, 1, 8, 0, 42, 10, 5, 26, 8, 1, 14, 29, -31, -2, 13, -41, -17, 0, 44, -25, -8, -1, 5, -9, 19, 11, 0, 25, -6, -11, -20, -41, -19, 21, 39, -8, -33, 16, -31, -14, 42, 6, -8, 13, -18, -25, 2, -4, -7, -5, 15, 19, -6, 9, 22, -41, -5),
    (-12, 14, -19, 3, 13, -2, -25, 8, -29, -25, -8, 13, 26, 12, -31, -5, -12, -6, -9, 8, 10, -2, -49, 10, -6, -14, -3, -9, 23, 6, -41, 16, -1, 1, -30, 13, 7, -3, -33, 7, -18, -10, 13, -8, 16, 15, -4, -9, 12, -21, -30, 5, 11, -11, -23, 14, -16, -9, 19, 22, 12, -22, -40, 17, -11, -11, -16, 10, 16, -35, -16, -19, 6, -17, 25, -9, 47, -5, -28, 8, -14, 4, -25, 8, 4, -8, -38, -2, -28, 16, 13, -8, 33, 8, -18, -3, 16, -23, 6, 2, 12, -14, -8, 8, -8, -4, 14, 0, 15, 9, -8, -22, 15, 4, 18, 2, 28, -27, -44, -9, 3, 14, 16, -28, 26, -9, -38, -22, 14, -9, -11, 13, 0, -11, -27, -25, -16, 5, 4, 1, 17, 3, -12, 0, -3),
    (-16, 16, -40, -6, 19, 28, -10, 30, -43, 1, -14, 26, 4, -7, -31, 24, 5, -2, -2, -29, -3, 17, 11, 24, 1, 27, -14, 2, -26, 0, -24, 0, 28, -23, 14, -15, -21, -8, 28, -5, 23, -31, -7, 7, -25, 6, 28, 8, -24, 0, -16, -18, 20, 41, -24, 31, -35, 4, -11, 17, -6, -28, -30, 16, -13, -2, 9, -30, 20, 1, -15, 29, -14, 8, -6, -11, -33, -30, -10, 12, 12, -8, 2, -22, -21, -2, 24, 2, 35, -23, 9, -15, 3, -12, 18, -14, -22, 0, -10, -26, -1, 37, -35, 21, -39, 30, -12, -12, 2, -36, -35, 17, -5, 1, 26, -17, 18, 8, -11, 17, 13, 6, -14, -22, -15, -20, 15, 6, 6, 17, 2, -10, -17, -1, 9, -7, 26, -1, -10, -18, -6, 3, -1, -10, 2),
    (-31, -31, 38, -36, -10, -11, -22, 13, -29, 15, 9, -13, 3, -47, -13, 16, -28, -57, 20, -1, 4, -22, -5, -13, -9, -20, 24, -20, 17, -31, 29, 1, -27, -2, -15, 8, 10, 7, -13, -18, 10, 25, 19, 2, -15, -12, 28, -27, -30, -59, 54, -54, 3, 28, -4, 4, -25, 31, 7, -1, 8, -59, 22, 20, -27, -24, 20, -40, -14, -12, 22, -3, -29, -25, 12, -16, 5, -45, 8, 1, -14, -6, 2, 15, -16, 28, 24, -12, 8, 4, 1, -11, -3, -47, -15, -11, -32, -43, 28, -21, -1, 49, -24, 6, -32, 2, -2, 15, 4, -51, -18, 46, -19, -25, 37, -23, -8, 12, 7, 5, -9, 5, 10, -8, -15, -22, 17, 19, 12, 6, 19, 0, 1, -1, -9, -14, -3, -25, 6, 2, 12, 5, 13, -1, -1),
    (20, 34, -10, 29, 0, -4, 22, 16, -25, 25, 18, 14, 31, 27, -14, 8, 14, 28, -27, 33, 1, -1, 15, 23, -24, 18, 13, -26, 37, 25, 5, -15, -9, 6, 1, 5, -13, 20, 5, 19, -17, 1, -1, -39, -5, 15, -1, -22, 26, 11, 5, 41, -3, -23, 34, 5, 9, -9, 30, 16, 22, 13, -10, 19, 0, 5, 1, 30, -9, -23, 3, -2, -21, -1, 47, 7, 32, 6, -20, -20, -7, -11, -20, -6, -28, -35, 19, 15, 14, -9, 18, -8, 8, 4, 26, -2, 11, -9, 0, 27, -15, -54, 11, -11, 0, 3, 23, -13, -5, 20, 12, 1, 3, -13, -16, 14, -23, -26, 18, -16, 5, -25, 27, -7, 8, 19, 16, -24, 12, -7, -18, -16, -28, -43, 27, -4, 14, 2, -3, -32, -25, 6, 33, 2, 8),
    (-5, -3, 10, -4, -23, -19, 9, -9, 4, 31, 4, 24, -5, 6, 6, -7, -6, -16, 1, 19, -12, -18, 17, -11, 11, 17, 21, 2, 12, 7, -5, 17, -13, -16, -32, 9, -10, 9, -17, -4, -9, 25, 9, 22, 10, -16, 0, -8, 3, 9, 5, 10, 9, -25, 1, -21, -8, 21, -9, 6, -5, -5, -5, -5, -33, -22, 26, -10, -12, -33, 17, -16, -27, 22, 19, 16, 8, -24, 6, 8, -17, -3, -15, 3, 8, -8, -42, -8, -27, 25, 8, 5, 5, -14, -44, 22, -10, 14, -34, 2, -26, 13, 3, 8, 8, 9, -39, 13, -29, 3, -3, -3, -28, -13, 11, -16, -8, -7, -29, -2, 2, 22, -2, 11, 15, -23, 7, -13, -7, -12, 8, -2, -6, -6, 7, 0, -8, 32, -3, 8, -2, -19, -34, -4, 0),
    (-22, -20, 15, -24, -27, -9, 7, 21, -3, -3, -9, -17, -25, -3, -12, 1, 22, -28, 27, -4, -37, -13, 29, 5, 39, 26, 28, -12, 4, 32, 13, -11, 10, -18, 24, 20, -19, -3, -7, -2, 34, -6, 11, 20, -49, -9, -5, -26, -29, -42, -14, -24, -16, 33, -2, 21, 2, 3, -36, 9, -41, -3, -6, 14, 24, -22, 9, -25, -11, 8, -7, 14, -13, 18, 4, 0, -14, -11, 16, -4, -4, -13, -3, 12, -34, -5, 11, -17, 2, 2, 3, -31, -22, -10, 13, 20, 9, -9, -3, -1, 10, 15, -13, 23, 2, -2, -13, 10, -22, 5, -3, 13, 0, -19, -12, 0, 2, -15, -4, 4, -12, 17, -43, -5, -13, -18, -22, -38, -16, -24, -3, -32, -13, -5, 17, 34, 6, -20, -4, 17, -5, -13, 0, -15, -1),
    (-20, -27, 45, -2, -6, 0, -3, -8, -13, -17, 4, -16, -7, -30, -20, -23, 16, 21, -10, 6, 4, -3, -6, -8, 25, 6, 3, 6, -8, 5, -6, 19, 31, 38, -22, 13, 26, 1, 5, -1, -16, 16, -15, 21, 3, 24, 22, -10, -3, 3, 36, 41, -16, -23, -36, -13, -14, 9, 28, -15, 0, -6, 20, -18, 50, 13, 21, 37, -12, -48, -25, -13, 1, 19, 42, -10, 3, 26, 30, -24, 24, 20, 8, 28, 20, -24, -1, -21, 33, -11, 3, 7, -2, 26, 1, 5, -9, -7, 9, 17, -3, -3, -24, -15, -23, -8, 6, -23, 6, 12, 8, 9, 2, 6, -4, 18, -5, -32, -18, -34, 5, -3, 13, -8, 19, 45, 36, -3, -4, 1, -2, -9, -2, -13, 30, -13, 46, -10, 11, -23, 5, 23, 61, -5, -1),
    (3, -2, -12, -6, 21, -6, 3, 16, 21, 16, -2, 10, 29, 8, -8, 3, 3, -5, 8, -24, 36, -4, 13, 5, -3, -22, -9, 11, 15, 3, 17, -22, -16, 4, -9, -19, 5, -17, -2, -5, -33, -9, -3, 25, 12, -10, -3, 11, -9, 14, -14, -4, 29, -33, 10, 1, 22, 12, -38, -10, 3, 8, 23, -2, 4, -21, -27, -37, 39, -30, -8, 4, 30, -1, -9, -7, 9, -10, 21, -19, -2, -10, 15, -6, 10, 5, 1, -15, -17, -7, -15, 7, 32, -23, -21, 16, 18, 12, 3, -11, 20, -16, 30, 24, -3, -17, -37, 7, 4, 10, 46, -4, 14, 3, -18, -25, -1, -2, -5, 13, 11, -22, -33, 20, 28, -21, -17, -13, 0, 10, -27, -11, 13, 2, -19, -2, -6, -5, -19, 19, 16, -14, -32, 12, -3),
    (-24, -4, -8, 20, 13, -14, -7, -12, -9, -9, 46, 2, 17, 4, 12, 13, -10, -18, 9, 8, 3, 1, -3, -10, -27, -12, 43, 21, 7, -1, 0, 8, 17, 2, -26, 32, 7, 5, -6, 6, -23, -9, 8, 10, -2, 3, 3, -5, 3, -12, 27, -2, -24, -33, -13, -42, 20, 12, 38, -25, 34, 11, 24, -10, -39, -17, 20, 20, -41, -34, -17, -45, 1, -22, 34, -7, 2, 9, -10, 20, -27, -48, -5, -12, -36, -44, 5, -8, -1, -3, 32, 5, -26, 17, 11, 0, 21, -6, 23, 9, -12, -10, -16, 5, -20, 26, 16, -3, 17, -16, 0, 23, -11, -28, 30, -9, 12, -25, 2, -14, 15, 5, 23, 11, -18, -29, 26, 21, -31, -37, 10, -32, -20, -11, -10, -28, 8, -12, 10, 0, -2, -23, -4, 21, 3),
    (27, 16, 31, -8, -15, 5, -8, 13, -1, -30, -29, 7, 7, 24, 22, -37, 26, 20, 18, 25, 2, -3, -5, 16, -10, -13, -5, 9, 23, 6, 15, -23, 23, -3, 0, 25, -24, -23, -16, 4, -18, 1, 24, -11, 37, -7, -10, -19, 7, -39, 22, -4, -19, 38, -24, 22, -10, -27, 35, 14, -22, -8, 15, 5, 15, 8, 30, 13, -8, -5, -38, -14, -31, 3, 9, -2, -7, -6, -15, 7, 14, 12, 8, 14, 16, -25, -15, -19, 11, 17, 29, -5, 19, 8, -1, -1, 0, -41, 16, 3, -40, 6, -14, 21, -13, -9, 40, 0, -10, -44, 2, -13, -5, -44, 19, 17, 0, -17, 16, -28, 13, 18, 44, -9, -23, -35, 10, -30, 2, -11, -38, 18, 22, -17, 7, -40, 13, -4, 15, 1, 22, -20, 11, 11, 6),
    (9, 13, -26, -15, 0, -21, -33, 27, 0, 11, 2, 5, 10, -20, -6, 2, -3, -2, 3, -10, 16, -3, -5, -14, 5, -17, 1, 17, 16, 7, 41, -8, 3, 11, 28, -9, 12, 7, 32, 8, -12, -6, -11, 16, -10, -12, 30, -3, -11, 2, -3, 8, -8, -16, -3, 17, 7, 32, -2, 7, -1, -11, -6, -1, -12, 9, 17, -6, -9, 4, 26, 3, -2, -1, -10, 16, -10, -3, -5, 16, -7, 13, -2, -8, -21, 13, 36, 1, 15, 25, -37, 23, -14, -7, -10, 5, -6, -5, 18, -12, 27, -36, -1, 21, -18, 35, 35, 22, 10, -27, -37, 31, 4, 17, 15, 24, -11, -22, 20, 5, 25, 13, -5, 0, 0, 3, 6, 38, -9, -4, -17, -2, -4, -5, 19, -1, 11, -10, -25, 17, 19, 25, -3, 20, 1),
    (5, 13, 2, 5, 7, -12, 2, 12, -31, -9, -8, -23, 11, -7, -21, 8, -2, 13, 16, -10, 17, -8, 9, 14, 4, -3, 2, -6, -10, 12, 9, 19, -17, 8, -19, -15, 18, 10, 15, -14, -13, 8, 0, 6, 19, -20, -23, 11, 15, -17, -7, 2, 31, -24, -7, 9, -15, 4, 0, 22, 12, -4, 11, -16, 3, 1, 4, 4, 24, -10, -39, -13, 11, -13, 8, 22, 25, 6, -16, 13, 1, 15, -28, 7, 9, 20, -12, -15, -17, -1, -3, 14, 30, 3, 2, -10, 10, -6, -5, -6, 4, 5, 13, -10, -13, -25, -5, -8, -1, 4, 4, -2, 6, 5, 37, -1, 13, -4, 16, -30, 3, -19, 2, 19, 22, -3, -29, -9, 10, 26, -11, 15, 6, 7, -25, -22, -34, -9, 12, 12, 34, -5, -1, -9, -1),
    (0, 13, -17, -15, -8, 22, -1, -14, -10, 7, -8, -32, -3, 18, -12, -24, 10, 23, -6, 21, -9, 4, 16, 42, 27, -13, -15, -10, 22, 30, 16, 1, 25, 32, -25, 10, -2, 7, -6, 34, -18, -9, -3, -3, 10, 5, 25, -24, 5, 7, -20, -9, -32, 38, 6, -16, -9, -3, -11, -16, -12, -11, -5, -5, 15, 13, -7, 18, -14, 11, -9, 15, 5, 21, -3, -12, 18, 41, 3, -21, 10, 42, -51, 14, 24, 4, -17, 15, -15, 18, -1, 13, 15, 36, -3, -28, 11, 14, 20, 19, -24, -22, -8, -60, -26, -22, 27, -31, -3, 28, 13, -17, -1, 6, 4, 18, -8, -25, 6, -18, -7, 7, 38, -11, -4, 41, -5, -28, -16, 1, 2, 15, 4, -6, 1, -7, -9, -15, 19, -17, -5, 14, 25, -15, 3),
    (11, -12, 3, -40, -37, 32, -5, -48, 27, 16, -23, 14, -45, -15, 20, -12, -5, 0, 25, -32, -5, 0, 9, -23, 28, -14, -53, -7, 0, -11, -17, -7, -2, 3, -46, 19, 23, 15, -28, -1, -8, -10, -14, 3, 7, 39, 0, -3, 8, 8, -9, 27, -22, -36, 15, -24, 7, 5, 1, -25, -17, -14, 6, 6, 38, 15, 9, 32, 3, -57, -4, -30, -4, -11, 13, 0, -18, 45, 20, -5, 14, 6, 1, -26, -19, -20, 1, -34, 8, 20, 27, -4, -15, 29, -5, 3, 42, -20, 1, 30, 14, -8, 22, -16, -24, -11, 19, 4, 26, 29, 6, -9, 22, -9, 9, 27, 3, -22, -28, -32, 17, 4, 14, 3, 28, -9, -6, -4, 1, 20, 6, -8, 6, -17, 9, -32, -11, -12, 15, -12, 36, -34, -2, 0, 5),
    (-4, 2, -9, -29, 0, -22, -28, 28, -36, 21, -15, 18, 9, 1, -22, -22, -7, 23, 3, -9, 20, -25, 5, 25, -24, 24, -21, 13, 3, 15, -14, -20, -13, 22, 0, 0, 12, 11, 38, -9, -30, 12, -7, 44, -1, 20, -22, -12, -14, -2, 0, -10, 7, 4, 34, 3, 13, 24, -8, -5, -5, -26, 13, 0, -23, 5, 2, -18, 8, -8, -11, 23, -22, 24, -21, 2, 15, -28, -9, -15, -9, 28, -30, -1, -2, -5, 9, 2, -14, 13, 6, 35, 30, 4, -4, 2, -31, 15, -24, -25, 12, 2, 11, 12, -20, 15, -11, 1, -5, -15, -24, 3, -22, 13, -9, -12, 15, 10, 4, 9, 1, 1, -14, 22, 5, -8, -1, -2, -14, 26, 8, 8, 17, 7, -3, -11, -38, -4, 4, -7, 18, -10, -17, -5, 1),
    (11, -24, -15, -4, -17, 21, 0, -10, 17, 6, 8, 24, -20, -5, -25, 7, -36, -31, -9, -27, -1, 20, -6, 5, -8, -15, 9, 21, 5, -12, -33, -11, -35, -15, -20, -12, 14, 28, -5, 6, -11, 17, 1, 20, 8, -13, -31, 16, -9, -37, 1, -2, -3, 17, -6, 5, 14, 17, 6, -1, -20, -14, 2, 23, -15, -20, -8, 6, -15, 12, -10, -7, -35, 2, 7, 8, 13, -33, -26, 18, -27, -25, 6, -8, -4, 18, -38, -14, -35, 13, 10, -3, 20, -11, -30, 2, -7, -24, 31, -6, -17, 14, 19, -12, -22, 16, 7, 17, -5, -3, -6, 0, -21, -30, 5, 6, 24, 2, -32, -15, -12, 5, 33, 11, -6, -22, -1, 10, -18, 1, 15, -4, -5, 14, -30, -29, -40, 0, 14, 17, 24, -8, -7, 15, 0),
    (13, -27, -20, 3, 3, 4, -10, 4, -20, 1, 4, 32, -16, -4, -40, 3, 19, -18, 21, 24, 20, -4, -21, -1, -31, 4, 16, 13, 0, 19, -16, 2, -12, -12, 5, -8, 2, -1, -45, 4, -37, 36, 1, 13, -20, 3, -36, -4, 8, -1, 8, 10, -6, -18, 11, 12, -10, -6, 21, 17, -35, -14, -24, -10, 50, 9, 26, -1, -13, -40, -11, 2, -14, 27, 10, 9, -11, 21, 9, -14, 0, 19, -16, 6, -12, 7, 16, 9, 13, 5, -26, 0, -26, 14, -30, -18, 18, 2, 18, 4, 4, -41, 26, -30, -16, -27, 15, -11, 31, 4, 6, -12, 3, 3, 19, 16, -14, -44, 12, -21, -10, -30, 12, -28, 8, 45, 12, 5, -3, -5, 13, -13, 2, -8, 31, -12, 12, -31, -1, -25, 8, 24, 0, 21, 0),
    (20, 32, -21, -3, 1, -10, 2, 25, -4, -13, -15, -6, -31, 13, 4, -32, 42, 34, 5, 21, -7, -25, 1, 17, 10, 8, -4, 4, -20, 11, 8, -24, 28, -13, 8, 22, -1, -1, -38, 12, 15, -5, -4, -12, -35, -6, -2, -15, 22, -17, -2, 20, 8, -22, -18, 2, -14, -27, 4, -3, 41, 25, -7, -14, 19, -2, 21, 38, 16, -28, 28, -10, 2, -11, 30, 5, 21, 9, -6, 14, -30, -8, 15, 4, 23, -12, -6, -8, 34, 13, 21, -1, 33, -7, 22, -25, 2, 12, -21, -10, 17, 0, -29, -19, -8, 7, -15, -1, 6, 2, -18, 33, -4, 3, -20, 6, 8, 0, -35, -29, -19, -13, 15, 8, 15, 19, 4, 0, -15, 4, -22, -6, -12, 24, -36, -16, -15, 5, 11, -16, 11, -8, 4, 34, -1),
    (-2, 6, -23, 24, 2, -8, 11, 15, -34, 6, -20, 5, -14, 40, 0, -8, 36, 18, -37, 19, 13, -46, 8, -2, 15, -2, -34, -7, 1, 54, 8, -33, -1, 31, 4, 19, 21, -24, -12, -3, -11, -18, -10, 18, -4, 48, -3, -18, 13, 30, -24, 24, -28, -5, 10, 22, 26, -34, -5, -10, 10, 76, 13, 6, -2, 27, 2, 2, 14, -24, 36, 7, 23, 15, 13, -28, 3, 31, 18, -20, 5, 23, 5, -20, -22, 17, 37, -33, 25, -12, 12, -18, 7, -16, 16, -2, -20, -25, -15, -9, -4, 18, -8, -26, 10, -2, -28, -4, 6, -11, 12, -24, -7, 4, -41, -3, 18, 13, -33, -3, 3, -17, -2, 3, -17, 8, 8, 2, 16, -1, -6, 12, -11, -4, -3, -15, -2, 28, 11, 24, -2, 27, 12, 16, 0)
  );
  ----------------
  CONSTANT Layer_4_Columns    : NATURAL := 16;
  CONSTANT Layer_4_Rows       : NATURAL := 16;
  CONSTANT Layer_4_Strides    : NATURAL := 2;
  CONSTANT Layer_4_Activation : Activation_T := relu;
  CONSTANT Layer_4_Padding    : Padding_T := same;
  CONSTANT Layer_4_Values     : NATURAL := 24;
  CONSTANT Layer_4_Filter_X   : NATURAL := 3;
  CONSTANT Layer_4_Filter_Y   : NATURAL := 3;
  CONSTANT Layer_4_Filters    : NATURAL := 32;
  CONSTANT Layer_4_Inputs     : NATURAL := 217;
  CONSTANT Layer_4_Out_Offset : INTEGER := 3;
  CONSTANT Layer_4_Offset     : INTEGER := 0;
  CONSTANT Layer_4 : CNN_Weights_T(0 to Layer_4_Filters-1, 0 to Layer_4_Inputs-1) :=
  (
    (6, -25, 17, -20, -2, 3, -35, -2, 3, -25, 5, 24, -29, -5, -4, -2, -19, 0, -3, -13, -11, 10, 1, 17, 11, -2, -19, -13, 0, -1, -23, -3, 9, -2, -8, -6, -23, -14, -7, -7, 8, 16, 13, -22, -31, 6, -14, 31, -8, 12, 25, 5, -2, 12, -48, -5, 0, -6, -32, 12, 2, -27, 3, 2, 19, 1, 21, 2, -16, 7, 6, 24, 24, 0, -21, 9, -14, -6, 1, -20, 5, -6, 6, -14, 5, 6, 6, -21, -19, 28, 0, 0, -1, 23, -23, -8, -20, -6, -5, -16, 9, 9, 27, -19, -3, -7, -3, 11, 3, 4, 20, 11, 8, 5, -12, 11, 7, -8, 3, 15, -12, 5, 27, 22, 5, -8, -13, -20, -2, -6, -19, 7, -19, 6, 20, -3, 26, -1, 8, 15, 7, -13, 26, 13, -15, -1, 1, -13, -13, 11, -10, -27, 2, 10, 23, -13, -10, -6, 12, -8, -12, 17, 6, -5, 18, -2, -18, -5, -50, -10, -10, -6, 6, 5, 0, 12, -6, -8, -4, 2, 15, -1, 36, -6, -14, 2, -6, 6, 18, -19, 9, -26, -20, -4, 22, 21, -10, -3, -8, 16, 8, -4, -11, -2, 6, -21, 25, -6, 17, -1, -15, 7, 17, -4, 0, 6, 1),
    (-8, 0, 14, 8, 10, 10, -21, -9, 26, 6, -17, 23, 15, 38, 43, 26, 22, 8, 2, -16, -6, 12, 2, 19, -14, -2, -5, 13, 8, -11, -19, 25, -1, -14, 7, 23, 5, 24, 26, -24, -12, 41, -10, 7, -10, 3, -5, 16, -10, 2, -32, -10, 6, -11, 13, 19, 7, -6, 5, 22, -7, -1, 13, 2, -27, 58, 20, -12, -20, -9, -21, -12, 16, 26, 4, 13, 8, 13, -7, -23, 34, 8, -6, 35, -8, 16, 16, 12, 13, 15, 12, -18, -24, 21, 20, 38, 20, 30, 13, -10, -5, -17, 6, -5, -5, -31, 16, 34, 2, 0, 36, 7, -21, 35, 11, -6, 2, -12, -3, -1, 0, 11, -23, -15, 10, -12, -6, 4, 7, -6, -5, 25, -17, -6, 16, -5, -12, 28, 17, -24, 10, -8, -8, -25, 22, 20, 15, 5, -16, 15, 0, -6, 13, 0, 28, 2, -9, 10, 2, 9, 9, 25, -4, -10, -8, 20, 28, 28, 5, 8, -13, -17, 2, 5, -23, -4, 6, -16, -8, 17, -9, -5, 39, -9, 8, -1, 7, -16, -8, -8, 7, -3, -16, -9, -6, 4, -9, -12, -22, 2, -2, -2, 17, 0, -13, -23, 6, 7, -9, 15, 3, -8, -5, -16, 3, -25, 3),
    (-3, -17, 5, 13, -22, 4, -4, -27, 13, 9, -13, -20, 18, 4, 1, 26, 17, 0, -15, -5, 8, -10, 15, 13, -15, -42, -5, 6, 2, 22, -9, -42, -3, -9, 6, -2, 8, -2, -17, -13, 9, 12, -8, -1, 16, 12, 12, -11, -20, -29, -13, 23, 2, 19, -16, -18, 7, 2, -15, -4, 10, -8, -8, 12, 0, 15, -8, 10, -9, 13, 13, -1, -14, -25, -9, 7, -11, -7, -11, -22, -10, 26, 8, -26, 7, -6, -28, 16, 1, 9, -10, 12, 8, 16, 5, -7, -36, -28, 19, 4, 16, 3, -32, -39, -2, 3, 9, -4, 26, 3, 6, 18, 12, 4, -7, -8, 15, 13, 25, -18, -15, -24, 29, 12, 16, -2, 0, -35, 0, 3, -13, -10, -15, 5, 5, 0, -10, 3, -12, 8, 6, -4, 22, -15, -12, -3, -6, 1, -4, 9, -14, 3, -5, 18, 2, -11, 13, 12, -12, 17, -12, -9, 12, 13, 8, -5, 15, -19, -17, -1, 16, 15, 1, -6, -29, -24, -11, 22, 4, 15, 21, -2, 7, 13, -11, 15, 25, -2, -12, 0, 28, -13, 1, -6, 17, 18, -14, 11, -12, -43, -5, -17, 9, 0, -11, -2, -24, -12, 9, 5, 36, -21, -3, -6, 13, -15, -5),
    (-35, 25, -2, 0, -4, 5, -42, -23, -19, -14, 20, 10, -22, 0, 16, -22, -3, -24, -4, -9, 4, 3, -23, 2, -35, 14, 8, -11, 14, 4, -26, 32, 8, 3, 33, -17, 5, -7, 7, 15, 6, -28, -32, -8, 8, 8, -17, 12, -21, -15, 0, -7, 3, 16, -7, 19, 15, 12, 25, 9, 18, 13, 17, 3, 27, -22, -29, 16, 19, 19, 4, 15, -11, -25, -18, 9, -15, 1, 9, 0, -27, -17, 14, -15, 15, -3, 34, -10, -17, 23, -30, -14, -14, 13, -4, -20, -20, -1, -8, -17, 5, -16, 20, 9, -6, -4, 7, -21, 7, -3, -20, 4, -19, -14, -7, -13, 11, 1, 3, -21, -32, 14, -14, -16, 18, -14, -4, -4, -12, 19, 14, 5, 7, -1, 2, 0, -11, -26, -33, 1, -12, 6, -7, -9, -13, -18, -29, 7, 13, 2, -11, 13, 19, 26, 6, 0, 4, 40, 39, 0, 17, 16, 27, -17, 26, 0, 7, -8, -14, -22, -18, 4, 2, -21, -32, 30, 28, -1, 12, 2, -27, 10, 7, -11, -15, -1, -1, -3, 10, 20, 6, -19, -5, -22, -4, -23, -8, 6, -19, -7, 21, -12, 21, -6, -18, -10, -5, -9, 5, 31, 10, 0, -5, -4, 5, -5, 3),
    (11, 5, -32, 1, -29, -21, -15, -7, -58, -17, -23, -3, -3, -8, -23, 4, -11, -2, 28, -1, -15, 2, -8, 2, 13, 10, -22, 9, -21, 23, 2, -19, -26, -2, -24, -21, -10, 0, -19, 11, 6, -27, 37, 4, -5, -33, 0, 3, -3, 20, -8, -2, 14, -3, -3, -11, -7, 13, -8, -16, 14, -4, 3, 18, 23, -21, 14, -2, 8, -35, 19, -5, 25, 4, -1, -6, 21, -9, 29, -8, 38, -6, -12, -7, -6, -7, -1, 10, -15, -16, 9, 13, 3, 11, 11, -6, 19, 7, 0, -24, 16, -7, 20, -16, 30, 21, -21, -14, 0, 40, 15, 20, 15, -14, -12, -8, -1, 22, 11, -3, 4, -25, -15, -19, -7, -10, -3, 16, 9, -10, -14, -7, 13, 12, -3, 6, 4, 22, -11, 12, -11, 8, -20, 2, 8, 17, 22, 1, 2, -9, 4, 2, -3, 8, 8, 9, 0, 16, -3, -14, -12, -13, 7, -10, -18, 2, 9, -14, -6, 25, -17, -18, 1, -24, -19, 19, -9, -12, -11, 14, 1, 18, 4, 13, 10, -30, 12, 0, -7, 22, 13, 12, -28, 9, -21, 11, -38, -9, -24, 11, 2, -20, 4, 1, -22, -1, -5, -7, 0, -28, 12, -4, -11, 31, -2, 5, 0),
    (11, 28, 20, 17, -27, 7, 26, 12, 8, 9, -5, 1, 0, -11, 26, 20, -12, 20, 18, 12, 0, -26, -2, 9, 0, 20, -15, -2, -25, -10, 47, 21, -15, 6, -8, -17, -5, -54, -12, -1, 8, 12, -3, 32, 8, -18, -17, 3, 7, -26, -10, -17, 0, 19, 24, -7, 21, 13, 3, -21, -17, -23, -40, -6, -22, -44, -23, 21, 16, 8, -15, -4, 17, 20, -20, 14, -11, 6, 19, -1, -14, -5, -1, -6, 0, -23, 5, 11, 3, 20, 14, -4, -11, -24, -6, 8, -3, -23, -13, 10, -13, -21, 44, 11, 6, 15, 11, -8, 2, -36, -14, -6, -9, 19, -7, 12, -5, -32, -34, -18, -29, -37, 11, -1, -1, 12, 25, -12, 38, -6, -2, -17, -27, -9, -33, 19, -8, -40, -34, -7, 1, 11, -15, -24, -5, -9, -2, 7, 4, 0, 7, 11, -1, -4, 28, -3, 4, -11, -4, -1, -2, 5, -10, -5, 11, -13, -16, -10, -28, 2, 14, 6, 9, 0, 1, -9, 15, -6, 13, -24, -24, -9, -12, -11, 9, 1, -15, 6, -4, -8, -27, -37, -25, -24, 9, -10, -3, 7, -7, -28, 52, -8, 6, -28, -19, 19, -19, -12, -13, -2, -4, 8, 8, 0, 5, -34, 4),
    (7, 10, -2, 11, -17, 13, -19, 4, -11, 1, -20, 9, 16, -19, 35, 19, -20, 12, 34, -13, 7, -1, -4, 9, 9, 8, -12, -4, -10, -5, 4, -25, -11, 6, 23, 21, 12, -9, 9, 15, -13, 46, 8, -15, -12, -12, 3, 9, 6, 6, 10, 14, -14, 10, 12, -1, -23, 1, 1, 25, -7, 8, -14, -8, 10, 20, 3, 7, -1, -27, -9, 11, 1, 18, 0, 5, 40, 15, -10, -9, 31, -2, -18, 4, -30, 22, 17, 3, 10, -19, 16, -23, 9, 7, 29, -5, 17, 27, 4, -8, 15, 11, 0, -19, 24, -3, -12, 24, -30, -6, -1, -12, 3, 10, 22, -29, 7, 20, 17, 12, 40, 31, 24, -6, -5, -2, -2, -39, 28, -13, -9, 25, -4, -18, -5, 1, -12, 30, 25, 2, -5, 3, 22, 18, -43, 7, -3, 9, 8, -1, -14, 22, 12, 1, -15, -8, -24, 21, 18, -5, -16, 8, -13, -3, -14, -24, 16, -21, -30, 21, 25, -19, -3, 2, -1, 11, 29, -15, -3, 16, -2, 21, -2, -21, -11, 31, 16, -21, -8, 6, 7, -9, -8, 5, 14, 18, -21, 11, -30, -25, 16, -20, -3, 8, -16, 5, -7, 13, 6, 7, -17, -2, -21, 0, 26, -1, -1),
    (22, 1, -2, 24, -20, 1, -11, -4, -36, -1, -17, 9, 30, 4, -13, 16, 4, -3, -1, 24, -9, 4, 6, 23, 15, 6, -17, 21, -32, 1, -26, 2, -70, -26, -10, 45, 1, -14, -21, 9, -9, -2, 0, 10, 5, -2, 6, 22, -18, -17, -30, 8, -13, 1, -6, -2, -56, -20, 22, 18, 10, -4, -22, -11, 15, -12, -18, -18, -11, -17, 8, 9, 19, 26, 1, 1, -1, 0, -6, -33, 7, -15, -24, -12, 1, 0, -8, 14, 3, -27, 11, 24, -13, -6, 22, 1, 27, 13, -13, 10, -2, 3, -14, -13, -15, -11, -21, -3, 19, -5, -20, 2, -12, -3, 15, 22, -3, 9, 23, 4, 0, 4, 3, 15, 19, -15, -6, -16, -18, -1, -10, 5, 30, -15, -12, 17, 25, 23, 8, -3, 22, 1, 2, 7, 20, -5, -5, -5, 2, 15, -4, -41, 9, -20, -5, -7, 3, -10, -19, -5, 3, -35, -11, 16, -4, -7, 6, -5, 21, -7, -1, 3, -4, 7, 0, -26, 3, 2, -13, -4, -8, 4, -41, -13, -16, -36, -29, 5, -11, -6, -1, 2, 5, -3, 9, -8, -2, 3, 13, -11, -3, 11, 8, -2, -7, -7, -20, 6, -17, -16, -30, 6, -27, 14, -15, 6, -4),
    (-1, 14, 16, 12, 21, 24, -2, -7, 0, 1, -12, 18, 5, 4, 37, 10, 6, -1, 31, -13, 15, 18, 8, 14, 5, -9, 4, 7, 10, 19, 22, -17, -5, -10, -10, 5, -15, 16, 7, -19, 13, 4, 13, -17, 8, 15, -9, -11, 11, -10, -10, -17, 8, -11, 13, -4, 15, -27, -18, -12, 6, 17, -34, 12, 14, 9, 3, -10, -14, 4, 7, -13, -39, -27, 16, 5, 13, 30, -23, -11, 0, -2, 9, -19, -4, 35, 26, 5, 18, -12, -17, -2, -6, -3, 26, -17, -30, -20, -12, -10, -9, -17, -23, 8, 0, 1, 11, -37, 3, 34, 8, -20, -27, -38, 5, 8, -5, 5, 3, -3, 0, 2, -14, 22, -11, 1, -15, -9, 6, 4, 11, -18, 8, 20, -42, -29, -6, -10, 31, -15, 13, 15, -4, 15, -2, -27, -14, -14, -9, 14, -4, 24, -32, 18, 12, 2, 10, -10, 0, -4, -7, -5, -2, 6, -11, 1, -17, -4, 11, -22, -26, -14, -10, -12, 5, 23, -21, 11, 18, -19, -4, -37, -14, -26, -10, -9, 10, 11, -10, -7, -18, -4, 28, 8, -7, 12, -12, 11, 2, -3, -13, -12, 2, 0, 5, -19, -41, 16, 17, -2, 32, -4, -8, -31, -9, 32, -1),
    (-27, -7, 11, -11, 23, -4, 0, 18, 2, 22, 17, -19, 2, 17, 12, -7, 15, 10, -19, 8, 5, 8, -22, -15, -13, -4, 8, -2, 19, 2, 3, 42, 18, 5, 22, -19, -5, 15, 1, -12, 23, -12, -12, 1, 2, 27, -15, 5, 4, 5, 9, -6, 7, 1, 1, 9, 21, 16, -5, 1, 6, 2, 9, 13, 10, -5, 6, 17, -3, 9, 13, 8, -28, -12, 18, -28, 8, -15, -41, 5, -32, -33, -11, 19, -12, 14, -16, -12, -18, -1, -9, -31, 0, 19, 18, 11, -19, -4, 21, -24, 13, -1, -5, 34, -23, -21, -3, 13, -29, 26, -35, -2, -3, -29, -17, 12, -16, 13, 22, 8, -2, -15, 4, -11, -7, -27, 13, 4, -36, -14, 6, 7, -16, -4, -24, -24, -8, -2, -16, -5, -23, 23, 2, 21, 2, -4, 12, 6, -2, 17, -6, 22, 10, 6, -6, -5, 19, 11, 9, 7, 18, -4, -7, -9, -7, -21, 9, -11, -6, 4, -9, -10, -4, 21, -8, 31, -8, 14, -5, -4, 0, 16, -1, 7, -14, 7, 5, -8, 24, 3, 9, -14, 5, -15, -34, 18, -29, 2, 23, 6, 5, 16, -1, -2, -3, 4, -22, 3, -12, 2, -8, 9, 12, 9, 5, -15, -1),
    (6, -11, 3, 13, -4, -13, -60, -10, -48, 8, 19, 4, -19, -40, -31, 5, -16, -7, 4, -28, -15, -32, -10, 5, -5, -7, 9, 6, -6, -11, -37, -28, -25, 1, 20, -24, -27, -25, -31, -8, -9, -13, 14, -12, 5, -23, 12, -15, -13, 4, -17, -13, -40, 11, -23, -27, -6, -10, 5, -30, -21, -15, -8, -13, -4, -30, 23, -34, -32, -14, 7, -15, 15, -4, -4, -5, -6, 15, -62, -37, -11, -8, 25, -8, -16, -15, 0, -1, 6, -4, 1, 8, -6, 15, 13, -8, 9, -4, 22, 4, 0, 10, -45, -40, 37, -6, 46, -19, 0, 7, -42, 6, 8, -27, 23, 18, 7, 18, -1, -10, 1, -7, 5, 9, -3, 12, -21, -27, 7, 6, 17, -15, -9, 4, -44, -18, 3, -15, 16, -18, -16, -19, -3, 4, -6, -14, 2, 16, 4, -2, -13, -29, 0, 5, 23, -13, 7, 3, -22, 5, -2, -10, -1, 5, -2, 8, 5, -12, 3, 17, -2, 15, 21, 1, -22, -32, 24, 5, 3, -16, -1, 23, -21, 18, 11, -25, 12, 10, 3, 22, 22, -12, 6, 12, 8, -11, -7, 14, -8, -21, 5, 2, -14, -20, 2, 8, 2, 4, 21, 6, 26, 18, 12, 4, 8, 6, 8),
    (22, -21, -13, -16, 6, -1, 2, -34, 20, -26, -25, -17, -17, -8, -6, -17, -4, 23, 18, 1, -22, 2, 5, 6, 13, -15, 13, 11, 1, 24, -11, -32, 11, -4, -6, 8, 15, -9, 14, -1, -1, 9, 4, 15, -25, -3, 20, 1, -3, -17, -6, 9, 9, -9, 24, 0, 1, 2, 1, 10, 17, 10, 12, -2, 10, -2, -11, 19, -4, 0, 1, -18, -1, -17, 1, -3, 19, -21, -26, -18, -20, -16, -23, 17, -20, -17, -3, -34, 18, 12, -18, -4, -25, 9, 19, 10, -8, -1, 35, 18, 2, 32, -32, -30, -15, -13, -6, 32, 14, -1, 22, 3, 8, 34, 13, -18, -14, -1, 12, 26, -10, -14, 1, 10, 6, 0, 6, 20, 7, 11, -9, 16, 9, -10, 26, -16, 8, 28, 6, 6, 14, -3, 5, -6, -35, -13, -10, -19, 5, 0, -37, -38, -11, -4, -12, 18, -14, 1, -10, -9, 8, 10, 12, 4, -2, -9, 15, -4, 10, 6, 13, 11, -1, 1, -36, -16, -5, -1, -17, 10, -5, -3, 10, -5, -3, 3, 12, 18, 17, 15, -2, 20, 4, 7, -16, 21, -7, -13, -1, -10, 0, -9, 3, 5, 12, -5, 17, 4, 12, 3, 14, 17, 15, -3, -1, -7, -2),
    (-29, -7, -28, 10, 6, -16, -9, -6, -16, -13, 3, 4, 8, -27, 28, 4, -15, 56, -20, -18, -5, -19, -9, -11, -18, -5, -34, 1, -18, 0, 17, -1, -12, -15, 0, -13, -12, -26, 15, 6, -18, 46, 4, -3, 10, -45, -31, -19, -3, -2, -14, 17, -33, -10, 19, 6, 8, 16, -11, -11, -7, -4, 9, 8, 5, 22, -7, -16, 10, -27, -3, -8, -10, 8, -37, -15, -16, 10, 0, -2, -15, -11, -3, -1, -16, -21, 12, -15, -9, 6, 14, 21, 3, -23, -15, -15, 13, -4, -41, 7, -41, -17, 31, -3, -6, -13, -19, -28, 14, -7, -21, 12, -4, 32, -14, -13, 13, -31, -21, -14, 17, -5, -18, 7, -37, -15, 11, 4, 17, -3, -25, -38, 2, -1, -19, 10, -2, 24, -22, 18, 16, -18, 2, -10, 6, 18, -19, 13, -33, -5, 19, 8, -10, -15, -8, 9, -3, -16, -6, 5, -7, 1, 13, 19, -3, -22, -12, -12, 23, 10, -38, 1, -40, -22, 22, 18, 15, 1, -6, -18, 6, -29, -29, 10, -1, -8, -23, -3, 3, 7, 0, -9, 14, -6, -15, 18, -27, -4, 10, 18, 22, 15, -11, -15, -9, -18, -21, 25, 19, 6, 6, 31, 8, 6, -8, 8, 2),
    (1, -26, -23, 14, -11, 8, 18, -1, 6, 1, -29, -35, -8, -17, -8, 8, -2, -9, -22, 9, -4, -4, 10, -16, 17, -23, 16, 26, -29, 12, -2, -27, 39, -13, -47, -48, 11, -20, -28, -6, -1, -6, -8, 18, -5, -2, 3, -1, 5, 10, 8, 14, -11, 1, -8, -1, 1, -32, -29, -10, 7, 3, -19, -12, 13, 4, -1, 10, -13, 2, -7, 9, -18, -39, -27, 18, 9, -4, -8, -6, 12, 9, 8, -28, 11, -17, -4, -4, 0, -28, -12, 1, 9, -3, -8, -44, -7, -24, 16, 37, 4, 8, -12, -50, 64, 8, -25, -28, 18, -6, -17, -9, 14, -24, -29, 5, 0, -5, -3, -19, 6, -18, 9, 29, 8, 10, 1, -24, 21, -18, -7, 6, -11, 2, -16, -22, 9, 5, -11, 2, -2, 9, 17, 6, -31, -33, 3, -9, 17, 11, -1, 12, -1, 13, 14, -23, 3, 7, 22, -19, 7, -9, -47, 14, 22, -9, -4, -38, -42, -23, 3, 9, 22, 30, -12, -21, 27, 4, 24, -14, -11, 11, 22, 10, 19, -23, -23, -6, -6, 12, -5, -17, -5, -14, 7, 16, 2, -7, 1, -8, 18, -7, 25, 15, 0, 4, 17, -5, -7, 4, -4, -11, 6, -3, 0, 9, 1),
    (20, 13, 15, 0, -3, 13, 14, 7, 23, -10, -12, -2, -8, -20, 11, -8, 5, -14, -7, -2, -13, 4, 13, 4, 41, 18, 24, -1, -16, 19, 18, -35, 7, -16, 9, 11, 13, -41, -7, 4, -24, 21, 19, -7, 1, -11, -6, 29, 40, 22, -15, 17, -23, -11, 10, -25, 13, -31, -13, 22, 10, -34, -14, -8, -6, 11, -13, -9, -23, -5, -9, 41, 23, 8, 16, 12, 18, -5, -12, -25, 23, -13, -4, -13, -7, -9, -5, -21, 9, -23, 5, -1, -18, 16, 18, 14, 32, 3, 3, 23, -2, 12, -1, -42, -6, -22, 11, -3, 21, -9, 7, -10, 18, -17, 12, -17, -14, 2, -13, 23, 16, -15, -23, 16, -48, -10, 5, -40, 17, 3, -5, 2, -1, -7, -28, -20, -9, -20, -23, 5, -27, 1, -26, 17, 17, -18, 16, 13, 2, 4, -9, -5, 5, -15, -34, 3, -3, -7, 13, -26, -3, -1, 4, -13, -17, 14, 3, 12, 12, -17, -1, -23, -10, 11, -5, -18, -19, 0, -13, 24, -4, -29, -24, 6, 12, 9, -14, -21, -2, 3, -20, 16, -24, -13, 0, -8, -33, -32, 1, -5, -23, -9, 2, -19, -17, -48, -21, 7, -9, -58, -44, -23, -31, -25, -34, -13, -1),
    (12, -8, -15, 5, 9, -12, 4, -19, -4, -32, 9, 28, -12, -26, 0, 1, -11, 6, -22, -21, -12, 24, -6, -14, 12, -33, -18, 15, -17, -6, 18, 9, -34, -29, -5, -19, 4, -10, 9, -2, -4, 27, -38, -14, 11, 13, -9, -15, 11, -6, -20, -15, -30, 4, 5, 20, -12, -14, -14, -16, 12, 3, 0, -18, -3, 1, -23, -23, 7, -9, -25, -14, -4, -14, 1, 15, 2, 18, -3, -14, 28, 2, -19, -6, 14, 1, 10, 14, 4, -12, -19, 7, 0, 15, 25, -2, -4, -40, -27, 30, -16, 4, -5, -12, 11, -2, -39, -14, 8, -31, 5, 11, -1, -5, -30, 0, 8, 15, -3, -2, -5, -31, -23, 27, -26, -13, 10, 5, 2, -3, -38, -2, 10, -19, -7, 0, 14, -8, -30, 5, -1, 12, -13, -4, -13, -9, 1, 3, 4, 2, 8, -14, 15, 17, -4, -17, 12, 20, 8, 25, -9, -20, 14, -1, -2, 22, 18, -8, -12, -35, 0, 15, 18, 18, -2, -22, 21, 22, -13, -22, -13, -3, 7, 13, 13, -18, 1, -7, 11, 11, 8, -16, -6, -13, -1, 17, 15, 5, -9, -8, 9, -2, -30, -5, 7, -13, 2, -1, 24, -2, 8, 5, 0, -2, 4, 5, -1),
    (-37, -19, 1, 4, 25, 11, -46, 0, -9, -4, 2, -2, 3, 2, 28, -17, 18, -28, -4, 2, 9, 2, 12, -16, -48, -8, 8, -24, 23, 5, -26, -5, -21, 15, 26, 0, -20, -10, 31, 3, 9, -34, -22, 5, 6, -7, 1, -7, -17, 0, 8, 0, 4, -7, -4, 15, 2, 28, -14, 9, -10, -26, 42, 16, 18, -24, -13, -3, -9, 2, -13, 2, -37, -5, 26, -5, 29, 27, -26, -2, 17, 26, 21, 3, -4, 9, 34, -13, 2, -11, 16, -5, 5, 9, 25, -8, -26, 20, 20, -4, 7, -8, -7, 1, -20, 9, 4, 11, -6, -23, 42, 10, 9, -23, 5, 4, 3, -18, -11, -9, -10, -5, -4, 8, 17, -21, 5, 8, 14, 28, 0, 10, -4, -24, 15, 14, 7, -11, -14, 4, -5, -16, -17, -8, -5, 4, 4, 1, -5, 13, -1, 11, 9, 5, -25, -14, -10, 21, 7, 15, 14, 1, -9, 20, -6, 7, 3, -2, -6, 17, 2, -2, -12, 1, 8, 4, 0, -8, -21, 1, -20, -11, 20, 9, 4, 2, 9, -5, 10, -16, 11, -17, 2, 1, -7, 7, -1, 6, 10, 2, 9, 12, -41, -4, -3, -15, -7, 23, -10, -3, 7, 14, -3, -20, -8, 5, -1),
    (-7, 11, -15, 2, -6, -13, 12, 40, -47, 5, 0, 10, -27, -17, -2, -9, -12, 9, -18, 10, -4, -53, -20, -18, -26, -20, -9, 17, -24, 28, 5, -14, 0, 15, -7, -28, -12, -28, 21, 11, -1, -6, -5, 21, 17, -36, 4, -22, -8, -26, 23, 6, 0, 19, -4, -32, 11, 12, -27, -14, 13, -12, 9, -7, 12, -12, -25, -2, 17, -1, 13, -14, -30, -13, -1, -5, 3, -3, -18, 27, -6, -12, 14, 7, -10, -5, 17, -7, 12, -14, -22, -9, 19, -45, -6, -31, -60, -38, -7, 26, 9, 28, 2, 17, 0, 25, 26, -30, -14, -26, 37, 10, 6, -28, -18, 13, 8, -36, -6, -46, -31, -11, 10, 0, 11, 28, 2, -7, 22, 1, 24, -7, 0, -21, 27, 9, 27, -32, -21, 9, -11, -16, -7, -18, -14, 11, 17, 6, 13, -8, -18, 12, 19, 19, 17, 7, -16, 1, -15, -4, 0, 9, 13, -9, -21, -18, -2, -4, -26, -7, 14, 16, 11, 10, 1, 16, -7, 1, 20, -6, 1, -16, 8, -5, -5, -3, 4, -5, 12, -17, -20, -23, -12, 6, 6, -4, 7, 7, 7, 6, -3, 13, 26, 8, 1, -9, 24, 7, -8, -1, -21, -11, 7, -9, -19, -13, 3),
    (-10, -15, -19, -5, -18, -14, -33, 3, -30, 16, 44, 8, 0, -22, -3, -17, 7, -5, -35, -5, -22, -3, -7, -12, -11, 7, -38, 2, -22, -14, -12, -10, -31, -11, 20, -8, 1, -19, -18, -11, -4, 11, 6, -8, 8, -30, -13, 2, 1, -8, -27, -16, -10, -9, 9, -5, -11, -1, 17, -7, -17, -9, -28, 9, 2, 14, -14, 17, -11, -23, -7, 9, 10, -2, -19, -19, -3, -8, 0, -12, -6, 8, -7, 10, -15, -28, -29, 5, -11, -1, 18, -20, -8, -7, -15, 5, 26, 1, -13, 7, -6, -3, 39, -8, 55, -7, -11, 7, -8, -41, -36, 20, 1, 16, 15, 2, -3, 16, 0, 23, 20, -3, -7, -14, -29, -10, 27, -20, 17, 9, -9, -7, -11, -10, -6, 11, -3, 4, 1, 5, -17, -10, -10, 13, 10, 4, -7, -4, 17, -8, 26, -29, 32, -2, 0, -6, 2, 8, -18, 5, -3, -11, -22, 9, 14, 16, 1, 17, 29, -20, 20, 4, 7, 7, 29, -28, 58, 15, -35, -18, -21, 6, -23, 6, -10, -6, -13, -16, 8, 19, 9, 8, 22, 0, 4, -20, -9, -13, 3, -33, 36, -10, 7, -13, -6, 19, -9, 16, -21, -10, 22, -11, -22, 11, 5, -5, 0),
    (-9, -29, 1, 0, 9, -5, 7, 5, 11, 16, 19, -17, 7, 7, 9, 4, 9, -17, -15, 16, 23, 3, 12, -8, -14, 2, 0, -6, 20, 7, -20, -19, 4, 7, 7, -5, 18, 17, 28, 17, 9, -27, -1, 26, 9, 20, 19, -2, 4, 12, -1, -5, 17, -2, -8, -28, 10, -10, 17, 18, -4, 1, 24, 2, 3, -13, 9, 5, -2, -3, -2, 7, -26, -43, 12, -17, 29, 24, -17, 23, 14, 26, 12, -3, 1, 30, 15, -9, 7, -23, 0, -10, 0, 13, 0, -17, -41, -9, -1, 11, 29, 5, -37, -6, -7, 1, 25, -4, 13, 36, 20, -2, 23, -21, 0, -9, -13, 14, 15, -13, -15, 17, -4, 9, 8, 1, -13, 1, 3, -8, 25, -2, 6, 11, 18, -11, 4, -9, 8, -12, -22, 0, 4, -8, -20, 24, 0, -4, 34, -10, -21, -3, 19, 4, -18, 16, -24, 8, 18, -21, -8, 23, -10, -6, -12, 5, -8, 6, -36, 22, -2, -19, 11, -3, -32, -22, 1, -13, 6, 13, -6, 22, 9, 0, -1, 22, -6, -18, -8, 28, 11, -11, -20, -18, 3, -23, 1, -12, -29, -15, 4, -23, 18, -24, -29, 5, -8, -17, -41, 0, 12, -26, -17, 6, -25, -10, 2),
    (5, 5, 9, 8, -14, 21, -20, -15, -1, 24, 22, -3, 6, 1, -17, -6, -13, 0, 26, -1, 6, 12, 0, 1, 2, 4, -3, 13, 0, 10, -40, -54, -8, 22, 11, -17, 19, 3, -27, 7, 6, 2, 7, 0, 10, 12, 12, 4, -10, 7, 15, 4, 5, 10, -24, -31, 1, -8, -12, -9, 3, -10, -15, 5, 5, -10, 3, 15, 2, 15, -5, 7, 14, -16, -8, 14, -18, -3, 0, -52, -8, -11, -17, -30, -1, -27, -8, 10, 7, 0, -33, 22, -14, -2, -21, 3, 0, -20, -11, 24, -16, 24, -22, -46, -11, 5, -14, -45, 16, -21, -44, -2, 15, -2, 0, 22, 15, -4, -2, 1, -17, 4, 8, 4, -10, -4, -27, -28, 8, 2, -15, -17, 24, -12, -32, -15, 17, -32, -1, 5, 6, -12, 1, -14, 3, -38, -21, -1, -12, -20, -8, -57, 10, -8, -2, -5, 10, -40, -14, -25, 0, -10, -44, 13, -26, -16, -29, -5, -6, -33, -5, -4, -11, 9, 5, -56, 9, -1, 0, -29, 8, -35, 0, 7, 3, 17, -45, 15, 4, -17, -27, -10, -17, -21, -1, 13, -3, -16, 2, -4, 17, 8, -10, -4, -10, -30, 2, 5, 18, 7, -29, -4, 1, -12, -20, -1, -2),
    (-3, 4, -44, 1, 14, -16, -14, -6, -40, -1, 0, -4, 3, -28, 15, -10, -5, -20, -7, -25, -17, -14, -9, -9, -13, 1, -38, -12, -12, -8, -12, 11, -48, 8, -10, 18, -7, -33, 2, 6, 9, 2, -6, -5, -2, -13, 3, 5, -8, 4, -24, 4, -11, -8, -7, 8, -20, -9, 12, -2, -3, 25, 30, 4, 3, -10, 3, -32, 20, 14, -6, -12, -7, -15, -35, -2, -13, 8, 0, -12, -42, -22, -9, -6, -6, -32, -4, 22, -6, -28, 7, 7, 8, -12, 4, -5, 5, -18, -17, -16, 2, 3, 23, 6, -21, -29, -19, -14, -13, -40, -1, -2, 14, -32, -16, 1, -13, -11, -2, 2, 3, -17, -26, -20, 6, -6, 3, 11, -11, -8, 1, -11, -19, -12, 6, 11, -2, -11, -6, 10, 2, 8, -2, -4, 13, 1, -23, 14, 23, 21, -11, -16, 24, -6, -26, -21, 5, -9, 10, 22, 11, -3, 4, -4, 17, 15, 22, -14, -3, -18, -9, 27, 20, 20, 5, -19, 11, 12, -1, -15, 14, -35, -10, 0, 10, 8, 15, 1, -9, 10, 12, -4, -13, -25, -32, 31, 5, 12, -2, -5, 3, -13, 0, 10, -4, -19, 4, 9, 18, -13, 18, 0, 22, -9, 6, 1, 4),
    (15, -32, -18, 0, -13, -16, -27, -18, -43, 7, 17, -12, -22, -11, -4, -13, -12, 23, 9, -15, -12, 1, -17, 10, 43, 16, -8, -25, -29, -8, 25, -11, 1, -16, -28, -3, -8, -18, -4, 11, 9, 12, 43, -1, -4, 17, -8, 26, 17, 37, 8, 6, -19, -10, 1, 15, -5, -10, -8, 21, 14, 16, 17, 7, 5, 13, 37, -19, -18, 13, -6, 20, 6, -4, 4, -22, 24, 1, -27, -13, -36, -21, 23, 17, -6, 6, 4, -8, -3, 12, 3, -32, 12, 2, -1, -11, 26, 17, 16, -21, 8, -20, -6, -3, 7, -6, -4, 29, -19, -1, 18, -6, -8, 24, 42, -20, 1, 25, -5, 21, 5, 22, 9, -2, 6, -12, -1, -4, -21, 2, -20, 32, -14, 18, 19, 1, -20, 20, 28, 0, -9, -1, 11, 25, 9, 5, 5, 2, 2, -4, -39, 0, 1, 1, 18, 6, -9, -3, -8, -12, -17, 23, 6, 2, -24, 26, 13, -9, -13, 5, 2, 3, 7, 13, -26, 5, -9, -2, -10, 28, 12, 18, -5, 7, 8, 23, 18, -21, -9, 21, 21, 12, 10, 24, 3, -6, 9, -7, -26, 8, 1, -3, 0, 22, 17, 14, 14, -7, 9, 23, 32, 10, 8, 11, 28, 11, 2),
    (6, 14, 10, 31, 8, 8, -3, -29, 8, -16, -5, 11, -3, 3, 6, 3, 6, -8, 12, 5, -14, -1, -8, 27, 0, 10, 31, 21, -12, -1, 7, 9, -19, -10, 10, 16, 24, -6, 10, -13, -2, 14, -7, 4, -14, -8, -11, 23, 1, -1, 21, -12, 5, 0, 9, 19, -15, 6, 15, 10, 8, -11, 7, 2, 3, 18, -19, 10, 11, -9, -13, -2, 16, 18, 29, 11, 9, 7, 8, -26, -10, -1, -23, -2, -2, -20, 15, 2, -7, -13, 1, -16, -18, 7, 10, 26, 17, 21, 39, 13, 7, 18, 16, 11, -34, -9, 6, 10, 11, -28, 17, 11, -5, 3, -6, -10, -18, -33, -1, 23, 17, 10, 23, -6, -4, -4, -2, 14, -17, 5, 3, -2, 1, -15, 12, 9, 8, -4, -6, 14, -18, -16, -15, -4, 7, 3, 10, -1, 17, -11, -6, -8, 3, -31, -22, 7, -11, 7, 12, -2, 11, -17, -13, 5, -1, 4, 15, 3, 27, 13, 4, 6, -5, 12, 14, -4, -15, -25, -15, 6, 11, -22, 5, -14, 9, -20, -25, -16, -18, -28, 20, -3, 13, 16, 0, 2, -11, -3, 6, -19, -6, -5, -21, -5, 10, -32, -5, 19, 7, 7, -14, 12, 2, -2, 0, -3, 0),
    (-7, 6, 19, 17, 1, 30, 5, 26, 7, -26, -13, 0, 5, 5, -4, -1, 6, 6, -6, 4, 10, 5, -13, -2, -7, 2, 14, -3, -6, -2, 8, 15, 1, -16, -15, 3, -10, 11, -17, -1, 15, 30, -35, -5, 18, -5, 8, -22, -1, -12, -2, 17, 11, 14, 21, 27, -24, -13, -46, 3, 0, 23, 1, -3, 0, 7, -21, -9, -3, 8, 3, -7, 4, -3, -4, 23, -22, 27, -11, -3, -6, 6, -22, -7, 19, 23, 7, -2, 12, -1, 2, 8, 14, 0, 2, -6, -14, -28, -6, 48, -6, 48, -11, -25, -20, -19, 9, 2, 4, 24, -13, -11, 5, 5, -15, 8, -10, 6, 4, -12, -18, -18, 14, 21, -5, 26, -10, 0, -11, -23, -13, -12, 2, 16, 24, -11, 13, 7, 3, 3, -10, -25, 16, -12, 4, -5, -22, -2, -28, -12, -6, -11, 10, 7, -19, -18, 14, -2, 17, 15, -10, -6, -26, -4, 18, 7, 6, -3, 0, -22, 8, 33, -11, 19, -8, -20, -18, -8, 18, -21, 18, 3, -21, -12, 10, -15, -4, 3, 11, -5, -3, -3, -8, -13, 3, 23, -7, 23, -6, 6, -22, -6, -36, -9, 12, 12, 9, -15, 24, 1, -19, 5, 3, 23, 13, 4, -5),
    (-2, -6, -14, -1, 15, -17, 7, 1, 34, -24, -25, 14, 0, 20, 26, 5, -16, 40, 25, -36, 8, 13, 9, 2, 21, -4, 7, 0, -15, -29, 16, 9, -17, -1, -10, -3, -6, 17, -8, 5, -5, 28, 5, -9, -9, 17, -3, 10, 28, -3, 3, -6, -15, -14, 18, 28, -25, 28, 1, 7, 2, 2, -17, 3, 2, 14, -10, 12, 11, -2, -3, 15, 20, 10, 2, 17, 6, -18, -18, -19, 40, -20, -11, 0, -22, 47, 13, -1, -24, 12, 25, -4, -16, 29, 12, 24, 14, -37, -29, -4, -2, -13, 25, -2, -35, -13, -6, -8, -21, 5, -17, 6, 6, 21, -2, 1, -8, 15, -18, -7, 21, -24, 6, -37, -15, -16, 23, 8, 16, 2, 1, 0, 14, 5, -14, 9, -16, 22, 4, 5, 6, 15, -24, -10, -20, -12, 3, -16, 0, 2, -16, -7, 37, -15, 12, 10, -12, 6, -5, -15, 10, 9, 19, -8, -10, -22, 5, 1, -4, -17, -8, -10, 12, -17, -5, -13, -14, 16, 3, 5, -14, 6, -38, -3, -21, 0, 11, -14, 1, 2, -7, -3, 27, -24, 3, -4, -3, -15, 11, 12, 19, -7, -4, 0, -9, 10, -31, -15, 0, -9, 3, -4, -4, 18, -29, 6, 0),
    (-7, 1, -10, -10, -14, -5, -21, -14, 3, 2, 29, -36, -20, 2, 22, -37, -13, 27, 5, 3, -5, 12, -4, 33, -13, 27, -7, 31, -25, 15, -32, -28, -2, 4, -5, -36, -13, 1, 0, 7, 5, 7, 22, -15, -19, -13, 3, -9, -7, 10, -14, -1, 5, -16, -1, -4, -19, -35, 10, -20, -21, 13, -7, -30, -27, -28, -24, -8, -21, -31, -4, -23, 6, -12, -17, -31, -3, 7, -37, 11, -48, -10, -28, 6, 16, -23, 12, -25, 13, 24, 10, -8, 10, 19, 0, -26, 12, 5, 21, -7, 1, 5, 18, -13, 30, 1, -28, 0, 23, -2, 14, 3, 3, 19, -2, 29, 4, 0, 0, -1, -2, -21, 1, 0, -8, -4, 7, -16, 13, -12, 5, -6, 13, 9, -9, 12, -8, 3, -3, 3, -10, -14, -3, -11, -34, -21, -14, -18, 2, -18, -30, 6, -18, -1, 10, 0, -22, 10, 2, -9, -26, 1, -17, -21, -4, 6, 2, -1, -19, -23, 28, -7, -14, -8, 0, -13, 7, -7, 26, -20, -6, -9, 17, -18, -23, -4, -5, -2, -8, 6, -21, 1, -15, -17, 0, 16, 7, 3, -24, -18, 28, -12, 1, -26, 2, 10, -7, -34, -22, 14, -10, 11, -29, -10, -17, -14, 0),
    (-13, 23, 2, -9, -1, 8, -31, 5, 8, 11, 10, 6, -12, 12, 15, -30, 11, 22, 1, -25, -15, 2, 10, 6, -24, 21, 27, -12, 13, 12, -20, 19, -11, -27, 5, 24, -6, 5, 44, -14, 12, 10, 25, -24, 1, 9, 16, 17, -5, -5, 4, -6, 8, 4, -2, 20, -11, 11, -19, 19, -6, -1, 35, 1, -12, 5, -5, -5, 18, 5, 1, 19, -40, 3, -10, 4, 16, -7, 13, 12, -9, 0, 6, 29, 11, 1, 20, -25, -13, 37, 25, -7, 6, 4, -9, 11, -11, 36, 23, 0, 7, -3, 11, 37, -14, -7, -17, 43, 5, -4, 49, -4, -12, 43, 31, 5, 7, 0, 25, 11, 4, 18, 1, 0, -2, -1, 11, 13, -12, 4, 2, 30, -7, -15, 45, 16, 2, 24, 16, -9, -6, -13, 17, 4, -24, -14, 5, -3, 32, -16, -19, -7, -13, -9, 13, 18, -14, 0, 27, -25, -18, 18, 3, -26, 19, -21, -15, 4, -6, 9, 4, -2, 17, 11, 11, 28, -9, 15, -27, 15, -18, -2, 37, 16, -5, 7, 13, -7, -4, 19, 9, 19, 5, 3, 4, -6, -12, -14, 9, 11, -13, 15, 0, 14, -2, -1, 15, 13, 1, 17, 14, -17, 13, -1, 2, 25, 2),
    (-16, 21, -8, -1, 18, -10, -50, -21, -51, -20, 16, 31, -13, 20, -8, -24, -17, 6, 10, -29, 8, -2, 7, -9, -28, -11, 1, 15, 8, 2, -6, -7, -18, -5, 36, 22, -20, 23, -20, -16, 3, 12, 16, -2, -12, -6, 9, -10, 7, -37, -7, -17, 27, -19, 2, 19, -8, -17, 17, 1, -19, -4, -20, -21, 0, 12, -29, -7, -17, 11, -2, -30, -16, 5, 10, 6, -7, 18, -43, -9, 17, 13, 18, 3, 13, 37, -10, -8, 0, -2, 34, 11, 5, 21, 13, -7, -25, 25, -6, -15, -2, 17, -40, -8, -7, 23, 33, 21, -1, 20, 1, -7, 7, 4, 24, -9, 22, 9, 15, 9, -18, 7, -26, -4, -2, -5, -4, 2, -9, 19, 28, -1, 8, 17, -6, -7, 0, -3, 19, 6, 10, 14, 7, -6, 8, 6, -2, 6, -7, -12, -2, -8, 19, 16, -18, -16, 22, 20, -9, 2, -15, -6, -5, -1, 18, 12, 15, -9, 3, 20, 17, 7, -10, 6, -12, -3, -7, 19, 14, -18, -8, 24, -11, -13, -3, 8, 29, 20, -6, 3, -2, -4, -2, 13, -3, 5, 0, 6, -19, 18, -29, 20, 0, -1, -4, 22, 3, 4, 0, 15, 4, -15, 5, 14, -1, 17, 2),
    (-18, 6, 0, 19, 7, 14, -7, 14, -16, 28, 18, -4, 12, 4, 11, 18, 3, 11, 20, 14, -10, -14, -3, 2, -20, 0, -30, 9, -16, -5, -8, 1, -30, 19, 19, -23, -7, -5, 22, -12, 17, 11, 19, 8, 10, -43, -1, -8, -14, -8, -38, -8, -42, -17, -7, -2, -11, -3, 5, -31, 6, -1, 17, -5, -24, -5, 3, -3, -2, -28, -18, -25, -33, 14, 8, 27, -4, 1, 15, 39, -23, 13, -14, 27, 4, 11, 30, 8, 25, 29, -2, -1, -11, -24, -6, -7, -40, 7, -4, 11, -4, 14, 8, 53, -49, 6, 8, 15, 22, -13, 61, 10, -7, 14, 8, 20, 26, -47, -9, -7, -16, -15, -34, -18, -26, -9, -7, 12, -16, 27, 23, -26, -11, -4, 1, -1, -3, -36, 0, 1, -10, -36, -2, -37, -17, 22, 2, 10, -15, 11, 20, 25, -15, -10, -2, 7, 13, 3, 32, -11, 7, 16, -17, 2, -11, -7, -1, -2, -28, -1, -2, 11, -7, 9, 6, 48, -18, 5, 7, 18, 17, -5, 49, -16, 16, 32, -20, -4, 5, -33, -13, -2, -21, -27, -9, 16, -1, -10, 3, 17, -4, 23, 33, -28, -15, -8, 15, -7, 8, -37, -23, -19, -7, -9, 2, -5, -1),
    (-7, -30, -3, 9, 5, 16, 10, 22, 13, 18, -39, 4, -16, 13, 1, 9, 16, -3, -17, -8, 13, 8, 9, 11, -11, -42, 5, 10, 21, 16, -12, 17, 9, -5, -28, 28, 14, 21, -8, -12, 18, -3, -29, -6, 16, 10, 9, 11, -6, -22, 0, -2, 8, 14, -2, 18, 3, 0, -23, 8, -13, 9, 11, 12, -5, 16, -12, -11, 17, 19, 3, 5, -19, -22, 16, -1, 17, 15, 5, 20, -6, 1, -31, 11, -2, 25, 21, 9, 18, -4, -16, -21, 32, 9, -13, 13, -18, -11, 21, -20, 30, 16, 1, 30, 14, 12, -4, 34, 8, 22, 42, 7, -14, -13, -19, -17, 26, 12, 4, 4, -5, -5, -13, -3, 15, 3, -6, 22, -7, -4, 5, 14, -4, 11, 33, 7, -1, 13, 4, 0, 2, -8, -3, 0, -6, -4, 27, -15, 5, -20, 5, 25, -11, 12, -19, 19, 0, 8, 34, -2, -24, 6, -11, -15, 8, 1, 6, 10, 9, 23, 6, -18, 20, -10, 14, 27, -28, 14, 17, 30, -14, 25, 37, 6, -8, 13, -3, -18, -5, -10, 10, 16, 14, 24, -1, -22, 2, -16, 8, 2, -20, -8, 32, 19, -2, -14, 24, 4, -8, 16, -2, 1, -13, -4, -8, 24, -6),
    (-4, -4, 11, 5, -5, 11, 5, 6, 11, 11, 10, 3, 5, 18, 8, -14, 1, 3, -1, -14, -6, -11, 3, -4, -34, -11, 27, -2, 13, 20, 3, 12, -25, -2, 41, 26, 16, 22, 41, 13, 9, 11, -42, 6, 27, -5, -5, -14, -11, -28, -24, -10, 13, -25, 20, 20, -7, 0, 18, 26, -11, 19, 7, -14, -27, 14, -44, 5, -5, -2, -32, -7, 2, -3, 19, 18, -4, -5, -9, -1, 0, -1, -1, 34, 22, 26, 35, 11, 19, 7, -23, -4, 0, 1, 20, 19, -7, 1, 15, 19, -11, 4, -7, 15, -16, -8, 51, 36, -6, 19, 21, 6, 20, 28, -8, -10, -17, -15, 2, 22, -2, -12, -24, -24, -5, -19, 32, 37, -25, -5, 10, 1, 6, 16, 1, -15, -13, -5, 9, -13, -9, -3, -20, -24, 13, -1, -4, 18, 1, 11, 2, 9, -7, -11, -18, 7, -8, 14, 12, 3, 5, -4, -20, 20, -23, 7, 4, 33, 34, 22, 9, 11, -51, 12, -1, 6, -8, 2, 17, -15, -10, -11, 22, -14, 5, 21, -12, -10, -33, 12, 17, 17, 6, 26, -28, -27, -22, -20, 9, -10, -4, 2, 30, -24, 5, 0, 13, -13, -7, 2, -6, 6, -5, -8, 10, -20, -5)
  );
  ----------------
  CONSTANT Layer_5_Columns    : NATURAL := 8;
  CONSTANT Layer_5_Rows       : NATURAL := 8;
  CONSTANT Layer_5_Strides    : NATURAL := 2;
  CONSTANT Layer_5_Activation : Activation_T := relu;
  CONSTANT Layer_5_Padding    : Padding_T := same;
  CONSTANT Layer_5_Values     : NATURAL := 32;
  CONSTANT Layer_5_Filter_X   : NATURAL := 3;
  CONSTANT Layer_5_Filter_Y   : NATURAL := 3;
  CONSTANT Layer_5_Filters    : NATURAL := 48;
  CONSTANT Layer_5_Inputs     : NATURAL := 289;
  CONSTANT Layer_5_Out_Offset : INTEGER := 3;
  CONSTANT Layer_5_Offset     : INTEGER := -1;
  CONSTANT Layer_5 : CNN_Weights_T(0 to Layer_5_Filters-1, 0 to Layer_5_Inputs-1) :=
  (
    (42, 2, 23, 21, -45, -14, -50, 3, -14, -18, 1, 2, 6, 35, -43, -24, 1, 14, -40, -52, -8, -41, -60, 35, -19, 29, 17, -30, -25, 41, 16, 39, 14, 7, 25, -31, -5, -28, -8, 1, 36, 20, -4, 16, -23, 34, -6, 1, 14, 21, -16, -61, 6, 6, -38, 38, 15, -11, 15, -30, -16, 24, 35, 71, 20, -6, -10, -73, 24, 8, 16, 11, 26, 7, -6, 13, -21, 14, -15, 39, 20, 11, 19, -27, -16, 14, -12, 22, 7, -29, 19, 14, 2, -11, 24, 29, 22, 15, 12, 31, -37, 15, 56, 25, -18, -47, -27, 45, -24, -30, 27, -24, 21, 16, 10, -33, -35, -27, -34, 0, -8, -52, 43, 1, -91, 16, 30, 26, 44, -15, -4, 12, -32, -3, 26, -26, -18, -42, -17, 49, -27, -35, 10, -24, 28, 17, -10, -45, -48, -32, -37, 34, 20, -49, 24, 28, -80, -8, 20, 36, 7, -16, 18, -17, -17, 8, -34, -23, -28, -21, 9, 33, -10, -8, -9, -48, 8, -8, -6, -47, -24, -52, 29, 20, -20, -15, 45, 41, -6, -5, 11, 9, -18, -23, -14, 1, 21, 4, 53, 27, 16, 40, -46, 21, -16, -46, 47, -14, 30, -38, 18, -39, -17, -15, -28, 26, -21, -62, 19, 19, -50, -6, 0, 10, -13, -30, 16, -5, 15, 13, 25, 4, 0, 7, -4, 24, -36, -79, 71, -11, 35, -31, 43, -97, -21, -21, 28, 34, -12, -61, 40, 37, -34, -1, 18, 22, 0, -14, -20, -36, -21, 31, 10, 8, -5, -33, -19, -4, 6, -31, 43, -68, 28, -26, 21, -79, -22, -18, 39, -20, 10, -19, 29, -2, -33, 8, -38, 19, -5),
    (-3, -39, -7, -6, 9, 10, 32, -1, 9, 22, 16, 33, 19, -2, -14, -10, 37, -32, -5, -28, 9, 21, 41, 50, -18, 23, -75, 42, 27, 54, -5, 3, 2, -81, -18, -30, -5, 76, -14, -28, -29, 14, -68, 17, 28, -46, -8, 14, 5, -71, -7, -46, 23, 18, -2, 37, -45, 39, -63, 37, -9, 78, -4, -32, -12, -4, 1, -9, 15, 48, 6, -21, 4, -10, -11, -4, 6, 2, -22, 6, -60, -27, -35, 35, -25, 4, -48, -10, -47, 9, -65, -25, 0, 17, 1, 9, 0, -9, -11, 8, 21, 4, 20, -30, -5, 36, -2, 19, 15, -20, -42, 10, -6, -15, -20, 25, -8, -18, 4, -31, -32, 49, 5, -9, 8, 31, 18, -18, -31, -33, -21, 39, -16, 27, 12, -54, -12, 1, -87, 5, 19, -7, -103, -27, 15, -35, -48, 42, 20, -27, -16, -61, -6, 48, -5, -21, -21, 47, 24, -51, 13, 10, 26, 11, -11, -35, 26, -27, 20, 7, -49, -22, -18, 43, -61, -24, -47, 17, -53, 84, 1, 7, 1, -43, 5, 9, -28, -32, -24, 12, -4, 14, -6, -43, 19, 17, -29, 30, 36, 7, 9, 36, 11, 28, -47, -21, -70, -21, -23, -11, -31, 23, 17, 0, 9, -23, 14, 14, -32, 6, -20, 24, 26, -2, -19, -5, 15, 53, -18, -19, -37, -30, 12, 42, -36, 6, -20, 28, -64, 0, 14, 30, -75, 46, 20, -9, -14, -40, -17, 23, -37, -14, 19, 10, 38, 2, -14, 20, 21, 10, -20, -58, 6, 12, 1, 7, -20, -5, -18, 56, 2, 23, -10, 29, -37, 22, 30, 9, 47, -15, 9, 47, 36, -16, -1, -1, 44, 9, 8),
    (1, 10, 26, 7, 26, -7, 8, -21, 28, 30, -36, 8, 36, -21, -7, -4, -14, 17, 4, 65, -26, 17, -1, -18, 27, -19, -47, 48, 34, -5, 12, 32, 19, 15, 18, -16, 23, 7, 9, -7, 12, 25, -10, 16, 31, -54, 13, 9, -28, 20, 28, 22, -67, -25, 3, -18, -2, 15, -14, 73, -22, -43, 16, 67, 35, 15, -34, -17, -19, 28, 15, 0, 27, 2, -30, 23, 9, -18, 45, -46, -5, 0, 25, 28, -22, -16, -5, 6, -33, 26, 36, 40, -27, -52, 29, 33, 36, 30, -24, -32, 29, -3, 37, -1, 30, 11, -42, 45, 9, -26, 32, -6, 2, 6, 30, 60, -14, -18, 23, -28, 18, -9, 46, 49, 25, 5, 26, 42, 16, 24, -22, 18, 28, -3, 35, -27, 52, 6, -33, 28, 36, -59, 30, 5, -7, 41, 44, 40, -37, -4, -30, -2, 12, -63, 47, 51, -21, 2, 1, 61, 37, 36, -18, -42, 29, -17, 14, -43, -3, 1, -6, -9, 13, 5, 53, 3, 44, 29, 63, 0, -37, -19, 22, -20, -27, -85, 34, 28, -31, -8, 41, 25, 8, -3, 7, -44, 16, -22, 29, 16, 50, 20, -12, 45, -29, -17, -10, 26, 22, -12, -21, -4, 19, -14, 13, 39, 9, 25, -5, 14, 13, 17, 28, 8, -8, 8, 3, 5, -6, -18, -6, -8, 8, 2, -11, 29, -34, -38, 2, -12, 34, 4, -21, 19, 10, 13, 21, 3, 16, -43, 52, -20, 13, -48, -19, 10, 6, -25, -5, -7, 2, 24, -13, -13, 32, 24, 9, -12, 7, 15, 1, 14, 26, 30, 27, 28, -22, 11, -2, -19, -20, -39, -26, 10, -14, -16, 4, 11, -7),
    (28, 14, 9, -19, -16, 24, 22, -29, 20, -8, 4, 33, 23, 27, -32, -16, 11, 9, 54, -7, 1, -36, -8, 26, 18, 12, -100, -32, -23, -20, 1, 43, -11, 47, -4, 8, 33, 3, 17, -9, 26, 1, -29, 33, -22, 6, -63, 5, -21, 20, 0, 31, 38, -45, -38, -9, -7, 12, -38, -36, -48, 3, -14, 55, 34, 29, -24, 31, 7, -25, -39, -49, 30, -26, 32, -15, 25, 1, 6, -16, -3, -16, -55, 24, 13, 23, 31, -27, 7, -49, 27, -44, 26, -8, 40, -1, -15, 52, 24, -5, 0, -20, 39, -26, -10, -43, -34, 34, 24, 17, -34, -64, -38, -9, 42, 23, 1, -1, 2, 13, 25, 30, -9, -32, -14, -23, -29, 75, 22, 58, 22, -13, 4, -51, 23, -18, 44, 12, -28, -5, -75, 15, -38, 7, -15, -10, -10, 52, 19, -78, 46, -2, -16, 24, 23, -26, -3, -3, -18, 51, 21, 58, -21, -18, -9, -11, -3, -5, 46, -29, 22, 22, 12, -21, -7, -29, -40, -55, -46, 15, -9, -33, 33, 23, 7, 62, -6, 2, -18, 3, 2, 23, 20, 43, 3, -15, 23, 1, 24, -22, 75, -16, 12, 32, 28, 40, -43, -5, -33, 15, -38, 18, 12, 3, -10, 21, 33, 9, -31, -8, 11, 1, -18, 23, 20, 18, 57, -34, 15, -22, -11, 18, 68, -6, 45, -3, -63, -1, -18, -31, -8, 1, -37, 19, 23, -21, 75, 13, 22, 13, -18, -15, 57, -5, -7, 48, -21, -11, 14, -16, 25, 23, 11, 16, 9, 27, -32, 9, -48, 9, -36, -44, 6, -67, -34, -5, -19, -9, 24, -17, -16, -4, -3, -43, 29, -6, 6, 27, -2),
    (-24, 2, 14, 17, -51, -3, -5, -48, 19, 21, 16, 2, 7, -17, -17, -4, -52, -39, -1, 44, 23, 33, 8, -43, -13, 39, 19, -21, 0, 63, 25, 25, 34, 11, -3, -1, -14, -42, -23, -1, 0, -8, 43, -10, 16, -35, -22, 48, -24, 3, 35, 33, 8, 12, 18, -47, -34, 49, -14, 20, 6, -12, 2, 41, 9, -13, -43, 49, 19, -14, -26, -17, 18, 1, 4, -35, 56, -24, -21, -3, -18, 28, 45, 23, -29, 44, -25, -50, 19, -16, 21, -3, -23, -32, -44, -29, -25, 4, -23, 57, -7, -39, 12, -32, 45, 34, 14, -19, 27, -28, 20, 33, -6, 14, 63, 32, 6, 41, 14, 8, -15, 54, 14, 2, 6, -7, 11, -43, -4, -15, 20, 15, 67, 25, -27, 4, -30, 38, 2, 12, -47, -6, 27, 35, 22, 8, 72, 32, -32, 45, -32, 13, -9, -12, 8, 38, 15, 68, -14, -31, -2, -50, -3, -7, 69, 52, 4, -17, -16, 16, 13, 6, 48, -3, 56, 31, 6, -27, 44, 10, 18, 47, -10, -3, -10, 12, 39, 34, 33, 52, 8, -34, -7, -33, -57, 40, -25, 16, 4, -13, -21, -9, -26, -11, 7, -11, 49, -22, -1, -49, 5, 53, -17, -48, -40, -24, -50, 40, 19, -5, -18, 51, 15, -38, -25, -22, -53, 35, -32, 33, 5, -23, -32, 10, -40, -16, 16, -26, 18, -75, -20, -20, 50, -18, -32, -25, -27, 2, -65, 43, 2, 10, -3, -9, -1, -27, 1, -6, -46, 15, -27, 9, -17, -10, -27, 14, -25, -46, -15, 4, 32, -50, -11, 37, 10, 36, -18, -41, -13, -17, 10, 0, 56, -7, 21, 3, 4, -27, 22),
    (24, 39, 5, 10, -28, 8, 1, -9, 10, -39, -33, 13, -42, -29, -3, -43, 49, -2, 4, 16, 16, 7, -4, -24, 21, -10, 15, 25, -23, 3, -30, 38, -1, 7, 11, 5, -55, 15, -42, -14, 7, -67, -13, 32, -5, 12, 7, -37, -4, 25, -20, 1, 11, 1, 22, 14, -8, 34, 6, -5, -51, 8, -32, 39, 12, -23, 30, 15, 16, -3, -27, 31, 20, -3, -7, 67, -50, -10, -1, -18, 21, -18, -23, -54, 12, -12, 65, 1, -1, -3, -3, 2, 14, 10, -11, 14, 13, -9, 2, 0, 11, -10, 33, -10, 29, 27, -3, -4, -25, -1, 2, -8, -9, -16, 14, 54, 1, 2, -8, 22, 4, 45, 46, -9, -11, 13, -25, 45, 79, 29, 42, -55, -11, 3, 21, -1, 36, -36, -32, 80, -44, -45, -75, -59, -20, 1, -45, 48, 18, -19, 36, 15, 4, 45, -6, 26, -38, 22, -6, 81, 43, 13, 40, -28, -27, 6, -25, -28, 10, -14, -1, 59, -16, -31, -41, -19, 1, -5, -28, 7, 24, -38, 37, -35, -27, -17, 50, 17, -4, 14, -34, 46, -40, -22, 2, -2, 13, -35, -20, 16, 39, 5, 11, 10, -17, 16, -48, -44, -45, -45, -19, 9, 39, 6, 5, 19, 0, 24, 28, -49, 9, 11, 2, -15, 67, -2, 56, -9, 8, -37, 31, 23, 43, 32, -13, 23, -43, -3, -39, -39, 4, -23, -28, 29, 6, 6, 15, 10, 28, 19, 14, -5, 11, 22, -7, 31, 5, -6, 23, 19, -10, 5, -21, -24, 9, -22, -2, 37, -31, -27, -53, -5, 8, -9, 2, -8, -18, -32, 28, 11, 29, -15, -17, 7, 10, 10, -36, 33, -4),
    (-30, 19, 28, -45, -16, 25, 7, 2, 3, -22, -44, -9, 31, 45, -30, 52, -1, 19, -38, 14, -11, -49, -40, -31, 26, 7, 24, -45, -67, -2, -22, 23, -39, 9, 1, 9, 22, 41, -4, -17, 9, 4, 46, -29, 41, 42, 9, 17, -33, 38, 0, 62, -13, 17, 40, -31, -6, -3, -3, -33, 14, -19, 23, 24, -20, 20, -30, 2, 51, 18, 46, 13, -15, 5, 46, -14, -13, 6, -3, -32, -34, -12, -21, 60, 16, 54, 12, -12, -43, 7, -35, -19, 73, -7, -3, 37, 11, 34, -10, 10, -10, -34, 26, 5, 30, 3, 35, 4, -15, 25, -46, -27, -55, -13, -4, 27, -14, -1, 67, -45, -23, 19, 4, -5, 20, -23, 54, -10, 18, 63, -17, 30, 45, -52, 11, -8, 54, 10, 21, 21, -51, -51, 40, -32, -6, -76, -18, 30, -38, 8, 29, -39, 0, 24, -52, 47, 23, -2, -3, 8, -13, 12, -27, 26, 1, -3, 6, -13, -4, 18, -47, 36, 0, -29, 59, 5, -10, -50, -47, -13, -14, -31, 25, 13, -7, -43, 11, 36, 9, 43, -42, 33, 26, 1, -45, -43, 30, -25, 31, -7, 50, 17, -22, 34, -52, -28, 78, -23, 22, -32, -18, -61, 21, 12, 15, -11, 7, 21, -3, 11, 26, -26, 10, 29, 22, -37, 9, -52, 47, -4, 18, 34, 9, 70, -12, 3, -36, -20, 22, 16, 9, 30, 0, -46, 14, 22, 46, 23, 31, 17, 19, 3, 0, 26, -15, 0, 5, -53, -7, -11, -13, 24, -13, 23, -32, 23, -4, -3, 9, -5, -2, 2, 24, 37, 25, 12, 17, 23, -37, 19, 28, -25, 7, 21, -37, 24, -17, -31, 8),
    (-18, -45, -17, 35, 7, -41, -9, -21, -21, 25, 39, -9, 33, -33, -21, 27, 15, 14, 27, 37, -15, 42, 8, -44, -22, 10, 45, 8, 20, 56, 27, -43, 9, -47, 12, 19, -6, -33, 5, -34, -12, -15, -4, 9, 35, 20, 32, 23, 28, 34, 34, 48, 17, 37, -48, 0, -12, -34, -13, -19, -43, 49, -1, -63, -6, -17, 21, 36, -13, -16, 27, -38, 4, 11, -19, -9, 50, 20, 41, 5, 20, 66, 56, 3, 7, 30, -46, -46, 7, -38, 39, 4, -6, 7, -7, -20, -13, -33, -26, -2, -40, 76, 9, 23, -37, 19, 7, 2, 24, -39, 9, 12, 29, -46, -12, -17, 17, -12, 53, -10, -13, -20, 19, 48, 35, 50, -26, -29, -34, -116, -22, 38, -54, 40, 12, -8, -64, 16, -31, -32, 26, -32, -2, 26, 30, -18, -26, -11, 21, -4, 61, 0, -5, 9, -26, 41, -11, 51, 2, -54, -39, -49, -8, 52, -30, -25, -30, -36, -62, -21, -27, -22, 19, -2, -22, 19, 13, -2, 27, -20, -23, 17, -23, -30, 8, 5, 14, 52, -28, 42, -11, -35, 6, -15, -25, -12, 12, 46, 20, -4, 43, 0, 3, 6, 2, 26, 28, 7, 19, -23, -9, -10, -9, -23, 29, 57, 9, -24, -30, 28, 27, 14, 2, 30, -17, -62, -8, 1, -30, 36, -21, 16, -18, 12, -16, -4, -2, -20, 8, 31, -5, -43, -11, -49, 7, -10, 18, 45, 1, -8, 43, 29, -17, 48, -39, 15, -51, -50, 10, 13, -21, -3, -43, -5, -33, -10, 1, -15, 13, -1, 1, 3, -16, 4, 7, 7, -4, -19, -39, 20, 32, 14, 18, 14, -58, 48, -46, 7, 4),
    (-68, 46, 37, 16, -1, -2, -8, -5, 19, -8, -56, -12, 2, -6, -35, 6, -49, -23, -4, 17, 32, -24, -45, 15, -1, 14, 23, -54, -10, -17, 12, -10, -9, 27, 10, 17, -10, -45, 35, 23, -14, 22, -50, -10, 30, 15, -38, 51, -65, -1, -30, 63, 15, -3, -73, 19, 15, 36, 42, -82, -60, -12, -3, 9, -4, 6, -21, 29, -3, -62, 29, 4, 1, -19, 10, 3, 7, 27, -9, 28, -44, 40, -14, 81, -14, 21, -35, -55, -20, 3, -34, -26, -42, 1, 10, -20, 8, -21, 10, 45, -5, -27, 14, 10, -34, 17, -46, -4, -42, 42, -24, 14, -16, -12, -4, 22, 26, -18, -31, 49, 18, -21, -29, -31, -50, -28, -2, 35, 19, -11, 54, 50, -65, -62, 6, 43, -43, 46, -11, 25, -52, 15, -92, 69, -6, 22, -42, 24, 18, 63, -44, 32, 1, 27, 68, -26, -49, -21, 59, 25, 27, 3, 38, 15, -52, -26, -25, 5, -14, 16, 17, 21, -30, 28, -73, 47, 22, 27, -31, 4, 26, 40, -27, 43, -26, 45, -2, -18, -35, 10, 34, 26, 15, -43, 25, 38, -27, -52, 51, 3, -45, -22, 2, 21, -37, 1, -21, 25, -35, -9, -9, -1, 2, 32, -16, 30, 14, 11, 31, 4, -38, 8, -15, 31, 36, -34, 12, 1, -36, -8, -7, 5, -39, 10, 18, 31, -36, -29, -37, 17, -9, 28, 4, -23, -18, 33, 14, -4, 7, 18, -15, 33, -22, 25, 13, 10, 31, -17, -9, -52, -23, 29, 7, -14, -5, -20, 1, 5, 2, 14, 8, 14, 18, 12, -10, -33, -38, -16, -17, 19, -45, 21, -40, 17, -13, -5, -19, -9, -8),
    (12, 41, -8, -19, -5, -24, -28, 37, 25, 12, -6, 34, -23, 11, -68, -22, 9, -12, -27, -20, 37, -21, 17, -1, 37, -5, 11, -26, 9, 66, -22, 33, 14, -21, 8, 53, 16, -37, 16, 2, 17, 36, 26, 40, -68, -69, -12, -51, 6, -40, -30, 8, 16, -36, 11, 21, 15, -37, 19, 16, 21, 32, -1, 39, 9, 13, 23, 55, -21, -10, 8, -7, -3, 8, -9, 34, -8, -61, 8, -19, -21, -11, -11, 3, -2, -12, -1, -4, -16, -28, 40, -54, 4, -5, -18, 29, -8, -21, -26, 0, -15, -8, 9, 26, 24, -4, -38, 30, 0, -2, -28, -16, -47, -30, 9, -12, 21, -22, 4, 25, 14, -12, -3, -13, -4, 51, -10, 50, -2, -20, 3, -12, 20, 15, 5, 51, -9, 26, -33, 64, -45, -34, -16, -47, -26, -80, 0, 11, 21, -39, 33, 29, 5, -30, 39, -21, 66, 21, -35, 35, -34, -27, 26, 35, -3, 23, 4, 17, -13, 11, -26, 9, -34, -69, -30, -14, -18, -25, -28, 1, 31, -34, 18, 10, -18, -55, 2, -16, -36, 13, -34, 15, 32, -27, -32, 17, 27, 19, 10, 4, 7, -6, 17, 37, -1, 7, 3, -6, -26, 0, 48, -8, 6, 38, -7, 11, -14, 18, 47, -1, -22, -8, -21, -28, 17, 14, 0, -15, 51, 15, 3, 37, 19, 17, 21, 54, -43, -34, -13, -19, -37, -52, -11, -32, 38, -20, 39, 13, 10, 5, -41, -30, 56, 38, -3, 1, 5, -7, 35, -18, -25, 43, -23, 8, -3, 8, -19, 6, 20, -35, -9, 25, -25, -18, -5, -36, 54, -38, -56, -3, 27, -38, -16, 2, -17, 17, -9, 19, -5),
    (-11, 49, 3, 16, -26, 12, -23, -14, -21, -54, 9, 17, 20, -1, -46, -83, -32, -15, -13, -22, 33, -64, -19, 4, -2, -38, 2, 3, -1, 32, -63, 43, -18, 16, -8, 24, 10, 11, -61, -14, -16, -54, 10, 3, 38, -1, -26, -57, -12, 13, -6, -6, 47, -39, -34, -24, 19, -31, 25, -34, -19, 17, 2, 21, -15, 5, -6, 7, 34, 3, -53, 9, 18, -32, 57, -10, -19, 14, -1, -17, -5, -9, -15, -36, 20, -10, 2, -14, 6, -17, -19, -19, -6, -20, 23, 3, 16, 0, -30, 12, 14, -20, 31, 5, 52, 11, 3, 0, 78, 32, -5, -20, -21, 56, 14, 86, 6, -12, -56, -27, -13, -44, 16, -10, -42, 3, -9, 32, 7, 91, 29, 23, 57, -20, 43, 20, 80, 20, -22, 8, 49, 15, -2, -49, -47, 42, -20, 102, 12, -25, -12, 11, -8, -2, 3, -45, -9, -8, 29, 58, -18, 54, -1, -16, 54, -33, 32, -8, 53, 15, 0, 2, 46, 1, 28, 3, -21, 6, -4, 23, -21, 12, 43, -16, -39, -4, 15, 23, 24, -37, -18, 28, -18, -67, 0, 10, 28, -25, -1, -8, -25, 13, 0, 27, -9, -14, -29, 23, -3, 7, -35, 46, -24, 13, -11, -33, 0, -4, -16, -49, 25, -19, -10, 12, -14, 23, -10, 33, 42, -48, 26, -9, 77, 13, 34, -9, -12, 1, 22, 6, 6, -2, -11, 54, -21, -23, -1, -10, -27, -37, 16, -69, 46, -34, -12, -1, 1, 54, 15, -13, -22, -19, 9, 9, 15, -35, 2, -45, 2, 3, 59, -4, 11, -40, 34, -6, 2, 30, 24, -29, -36, -31, -3, -45, 5, -18, -10, 6, 0),
    (-32, 5, -12, -15, -20, -22, -8, -29, -47, 4, -25, -25, 32, 4, -15, -6, -8, 26, -2, 24, -28, -41, -44, 16, -1, -16, -44, 38, -6, 18, -2, -28, -37, -14, -23, -28, -11, -11, 11, -6, -7, -20, -6, -39, 51, -6, 12, 14, 15, 9, 41, 31, -2, -17, -18, 18, -38, -14, 30, 58, 25, 27, 28, -29, -34, 14, -34, 10, 16, -8, -9, -25, 10, -20, 12, -15, 28, 0, 39, -31, 9, -4, 43, 31, -8, 0, 22, 25, 11, -16, 2, 44, 32, 5, -2, -12, -17, -37, 1, -19, 1, 12, 8, 24, -65, -15, -48, -10, 35, -1, 22, 78, -31, 17, 1, 34, -11, 51, -14, -27, 1, -28, -33, 51, -68, -6, 7, -20, -43, -12, -5, -30, 20, -15, 42, -4, -36, 1, -46, -47, 62, 9, 34, 72, -22, 32, 50, 27, -27, 38, -52, -11, -6, 1, -53, 38, -90, 12, 20, -21, -26, 20, -50, 11, 38, -24, -9, -6, 27, -10, 7, -11, 63, 2, 22, -19, -1, 1, 21, 18, -22, 6, -34, -47, -27, 12, -21, 1, -11, 26, 35, -15, -23, 19, 29, 6, 4, 16, 2, 8, 19, 19, -14, -30, 46, 8, 31, 56, -30, 41, 4, 19, -14, 23, -25, 3, -16, -48, 17, -5, -42, -16, 16, -21, -38, -3, 21, 3, 41, -5, 9, 17, 6, 46, -38, -36, 27, 48, 16, 70, -7, 43, 3, 20, 8, 56, -29, 23, 2, -4, -27, -18, -17, -27, 20, 12, 0, 7, 17, -3, 10, -37, 7, 4, 22, 4, -24, 3, 14, 42, -30, 22, 17, 39, -17, 18, -30, 39, -59, 8, 16, 3, -10, -48, -28, 0, 9, 36, -3),
    (-1, -22, -26, 32, -9, -37, 18, -17, 4, -1, 28, 23, -38, -5, -1, 8, -16, -28, -34, 8, 10, 26, 22, 28, 15, -35, -23, 26, 45, -3, 30, -46, 7, -30, 20, 11, -25, 25, 28, 9, 1, -18, 10, 18, -30, -59, 3, -6, -26, -4, -41, -42, 24, 7, 55, -34, 10, -12, -7, -9, 16, 67, 13, 6, -14, -22, 12, -2, -12, -36, 12, -53, -3, 14, 16, 2, 19, -16, 13, 13, -12, -22, 18, -47, -20, 8, 37, -23, 6, -2, -5, 58, -26, -24, -5, -1, -2, 14, 14, 4, 11, -18, 15, -4, 38, 30, 43, 20, -30, 30, 3, 7, 4, 2, -60, -8, 15, 37, 14, 4, -12, -2, 4, -16, 61, -35, -2, 34, -23, -10, -23, 23, 0, 65, -24, 16, 7, -1, 62, 4, -42, -48, 11, -5, 41, -32, -49, -78, 37, 15, 93, 4, -12, -20, 26, -26, 52, 11, 1, 6, -14, -41, 35, 9, -8, -3, -5, -22, -20, 23, 9, -21, -7, -29, -9, 36, 0, -2, 10, -34, 9, -12, 64, -36, 16, -57, 39, 18, -21, 2, 46, -48, -18, 19, -11, -15, 12, -29, 10, -44, 30, -1, -17, -9, -2, 28, 17, 32, -35, 19, 21, -2, -36, -11, -23, 13, 17, 14, -21, -22, -78, -30, 3, 13, 45, 3, -14, -54, -20, 56, -3, 12, 0, -28, 20, 3, 7, 19, 41, -21, -6, -17, 20, -33, 13, -36, -40, 34, -29, -16, 19, -18, -6, 23, -23, 8, -6, -15, -23, -48, -43, 0, -9, 28, -7, -57, 19, 2, -38, -10, -50, -28, 2, -26, -37, -48, 19, -7, -1, 33, -12, -45, 0, 10, 16, 49, -17, 24, -3),
    (-5, -2, -22, -37, -20, 32, 44, -7, -54, 13, -10, 40, -27, -16, 7, 5, -28, 7, 17, -50, 9, -9, 41, 23, 4, 36, -20, 24, -1, 37, -16, 44, -17, -41, 2, -2, -51, 18, 31, -5, -83, 10, -51, -8, 13, -19, -58, -40, -20, 42, -15, -71, 1, 0, -6, 27, 31, 15, 37, 33, -30, 20, 24, -17, 0, -43, 7, 13, -31, 17, 25, -2, -72, -7, -57, 29, -8, -13, -60, 20, 20, 26, -6, -1, -1, -31, 10, 7, 6, 2, -9, -6, -6, 13, 16, 17, -29, 11, 38, 3, -29, 21, 37, 8, -39, -1, -30, 34, -26, -38, -23, -9, -8, -2, -6, 13, -30, 14, 5, -4, -3, -13, 8, 2, -21, 36, 14, 14, -21, -31, 20, 58, -39, -35, 20, -5, -62, -10, -59, 15, -7, -35, 44, 15, 59, 60, 24, 16, -52, -29, 6, -6, -24, -62, 13, 54, -28, -3, 18, -2, -30, -18, -8, 40, -11, -37, 24, 11, -34, 21, -65, -5, -10, -14, 41, -11, 2, 80, 5, 6, -64, -16, -11, 16, -39, -38, 36, 30, -22, -5, 21, 32, -32, 4, 9, 13, -20, -31, 16, 15, -11, -6, -17, -1, -30, -36, 6, 4, 6, 14, -21, -16, -15, 42, 5, 16, -21, -20, -17, 7, -5, 27, 8, -37, 25, 8, 7, -8, 3, -37, 40, 9, -15, 16, 17, 9, -41, -38, 26, 34, 38, 6, 29, 41, -35, 28, -27, -1, -8, -69, -13, 21, 19, -37, -17, -7, 53, 14, 12, -3, 40, -33, 13, 12, 4, 6, 3, -16, -38, -23, 15, 41, -11, 32, 11, 7, -42, 3, 17, 25, -13, -40, 40, 33, -6, -58, 40, -51, 1),
    (28, -19, 13, -5, -16, -9, -8, 4, 3, -10, 7, -18, 3, 17, -12, -22, -6, 13, 10, 35, 40, -10, -5, 30, 39, -22, 30, -13, 16, 15, 1, 14, -34, 6, 50, 17, -49, 18, 0, 23, -39, 30, -20, -25, 12, -8, -5, 62, -6, 24, -68, 28, 39, 58, 13, 7, 18, 24, 9, 14, -22, -28, 26, 6, 1, 1, 14, -11, -18, 3, 18, 16, -38, 0, -18, -2, 7, 12, 22, 48, -9, -22, -2, 38, 26, 50, 32, 21, 32, 10, 50, 7, -60, -34, -25, 23, 0, -39, 6, -11, -16, 3, -7, 0, -25, 10, -10, -17, -20, -38, -10, -9, -2, -21, -15, -34, 11, -26, 31, -9, -47, 47, -63, -40, 28, -26, -19, -21, -8, -12, 45, -16, 1, -31, -54, 19, -20, 5, 28, -23, -50, 7, -37, 72, -2, 22, -14, -26, 35, 42, -3, -15, -23, 55, -10, -29, 57, -4, 19, -7, 26, -21, 20, 4, 11, -33, -6, 20, -1, 27, 50, 6, -29, 15, 11, 46, 48, 36, 8, 13, 2, 29, 0, 0, -23, -26, 13, -27, 26, -25, 16, -1, 8, -29, -46, 8, -4, -4, 1, -5, -4, -3, 43, 30, 55, -13, 26, 1, 11, -21, -7, -54, -32, 22, 12, -7, -2, 49, 9, 10, -18, 0, -13, -24, -6, -38, -57, -22, 0, -5, -10, -60, -38, -31, 26, -5, 39, -12, 40, 32, -12, -12, -12, -29, -20, 38, 27, -17, -5, 32, -22, -10, -29, 3, -34, -33, -26, -11, -33, -50, -3, 26, -35, -51, -58, -49, -10, -50, 21, 1, 42, -9, 43, -76, -10, 0, -18, 56, 10, -27, -43, 12, 22, 17, 14, 11, -27, -38, -6),
    (21, -3, 3, -31, -32, -31, -20, -13, 20, -20, 59, 25, -25, 21, 24, 9, 2, 45, 29, -13, -6, 38, -12, 10, -32, 10, -68, -45, 0, 9, 7, 6, 37, -15, -14, 6, -9, 28, 20, 9, 29, -7, 36, 41, 8, 15, 18, -43, 7, 42, 18, -52, -13, -23, -7, -14, -6, 7, -81, -10, 6, -15, 0, 36, -27, 28, -33, 12, 39, 51, -44, -12, -16, -4, 6, 26, 88, -29, -39, -13, 9, 17, 9, -39, -51, 2, -39, -29, -27, 16, -15, 8, -4, 10, 6, -18, 15, -37, -7, -32, 4, -28, 6, -28, 15, 1, 41, 6, 20, -24, 31, -17, 18, 32, 35, -65, -27, -2, -2, 0, -38, -39, -51, 26, 27, 30, 33, 0, 46, 40, -45, -35, 48, 62, 6, -2, 21, -26, 11, 2, 30, -49, 58, -53, 49, 25, 51, -59, -43, -47, -7, -23, -42, -12, -72, 53, 19, -11, -16, 10, -26, 4, -27, 27, 17, 64, -23, 9, 9, 14, 6, -3, 73, -4, 24, -31, 19, 6, 35, -19, -24, 9, -4, 5, -24, 8, -37, 5, 10, 4, -15, -10, 20, 9, -45, -11, 54, 31, -20, -26, 12, -5, -37, 26, 76, 13, 45, 16, 4, 26, 6, -30, -30, 28, -16, -18, -14, 33, -19, -9, -43, 5, -1, -45, -5, 8, -37, -40, 46, 35, -7, -27, -6, 11, -5, -26, 77, 15, 58, 8, 19, 32, 22, -5, -11, 10, -49, -31, 0, 4, -36, -6, -47, 3, 8, -67, -41, 11, -7, -2, 9, -22, 18, 9, 16, 21, -15, -7, 6, 24, 47, 21, 2, -10, 40, 0, 2, 1, -18, -40, -9, -1, 19, -3, 18, -32, 21, -2, -1),
    (-1, 14, -45, 13, -16, -18, -17, -13, -12, -33, 11, 22, -13, -16, -42, -7, -3, -32, 11, -37, -20, -15, -14, -32, -12, -20, 18, 11, -19, 8, -16, -37, 37, -8, 8, 10, -31, -23, 11, -26, -18, -52, -57, -3, 23, -43, -42, -9, -2, 1, 30, 27, -40, -21, -17, -35, 2, -57, -22, 19, -46, 35, -32, -8, 10, -3, -52, 41, -36, 11, -39, -19, -47, -84, -43, -10, 42, -32, -51, 21, -12, 46, 26, 24, -48, 28, -46, -23, -24, -69, 9, 43, -58, 23, -1, 11, 31, -34, -24, -12, 0, 27, -7, -18, 13, -36, 20, 10, 27, -72, -20, -47, 19, -16, 36, -45, -48, -29, 45, -3, -25, -10, 8, 57, -55, -2, -19, 4, 14, 2, -31, 19, 33, 44, 25, 1, 15, -31, -79, 41, 80, -6, 8, -49, 24, 0, 91, 1, -15, 4, 32, 13, -7, -6, -86, 20, -94, 19, 11, 11, -13, 52, 7, 66, 29, 1, 1, -9, 5, -22, -28, 10, 45, 4, 13, -14, 14, 16, 56, 76, -14, 0, -40, -53, -38, 14, 7, 39, -91, 31, -2, 26, 12, 17, -26, -23, 29, 64, 8, -3, 0, 13, -26, 24, 5, -6, 18, -9, 48, -15, 7, -10, -11, 24, 56, 6, -16, -25, -28, 55, -1, 38, 27, 14, 31, -19, -4, 1, 21, 49, 10, -8, 19, -5, -26, 2, 63, -29, -8, -6, 19, 5, 68, 11, -18, -17, 13, 13, -32, -10, -51, 41, -13, 34, 17, -9, -14, 28, 7, 41, 23, -10, -3, -40, 29, 16, -17, 1, 49, 14, 27, 10, -4, 19, 56, 29, -23, -36, -41, -2, -21, 26, -7, -9, -41, 7, 4, 17, 23),
    (11, 1, -49, 6, -37, -40, -5, -25, 9, 29, -14, 1, -54, 3, -57, -19, 10, -47, 1, 18, -44, -28, 31, 4, 15, 8, 17, 37, 18, 3, -41, 2, -12, 16, -13, 11, -13, 2, -48, -32, -22, 41, -32, 25, -19, -36, 1, -30, -3, -77, -55, 4, -31, -31, 18, 3, 18, -25, 77, 50, 32, 53, -31, 37, 9, 0, -55, 21, -31, 20, -44, 1, -1, 30, -31, -1, 34, -39, 24, 7, -39, -3, -24, 16, -11, -14, -21, -7, -17, 10, 73, -3, -58, 58, 5, -12, 18, -2, 18, 7, 8, 33, 6, 7, -41, 6, -11, 41, -49, -4, -24, -15, 6, 9, -1, -36, 13, -19, 28, 10, 12, -40, -28, 17, 36, 54, -5, 32, -16, 14, 5, 65, -17, -3, -18, -36, -21, -23, -72, 46, -1, -18, -5, -22, -22, 11, -43, 22, 17, -73, -14, 21, -3, -80, 7, 41, -23, 40, -59, 25, 7, 9, -1, -17, -35, -8, -31, 19, 29, -49, -4, -24, 27, 19, -14, 6, -8, -6, -13, 31, 1, -23, 26, 16, -3, -51, -35, 10, -58, -5, -27, -6, 29, -12, 16, -16, 7, 15, -11, 9, 7, 28, -1, 45, -13, 26, -45, 13, 29, 2, -3, 27, 3, -2, 20, 18, 44, -24, -1, -5, -17, 26, 3, 23, -42, -22, 36, 41, 9, 5, -18, -11, -20, 4, -61, -5, 10, 18, -42, 41, -34, 0, 23, 44, -7, -27, -40, 6, -27, -1, -4, -17, -28, 20, 10, 20, 41, 71, 8, -36, 38, -17, -23, -6, 20, -33, 22, 27, 21, 15, 40, -18, -17, 11, 32, -16, -19, -1, 13, 1, 4, 46, -9, 8, -36, -68, -19, 18, 2),
    (52, 31, 2, 0, 17, -42, -19, 5, 7, 12, 52, -11, -22, 31, -15, 25, 7, 13, 19, 4, -4, 26, 8, -26, 23, -3, -23, 32, 5, -58, -7, 1, 4, -1, 20, -23, 14, 7, -32, 7, -2, 19, 25, 5, -34, 4, -44, -12, 38, -19, 11, -58, 31, 39, 56, 4, -14, 45, -55, 30, 23, -25, -12, 3, 9, -33, -23, -52, 0, 50, -48, 4, -21, 4, 8, -4, -4, -5, -32, 10, 33, -13, -15, -59, 35, 25, 24, 23, -14, 38, -20, 3, -1, 18, 20, -10, 24, -14, -38, -27, 15, 35, -11, 10, -18, 1, 23, 10, -31, 22, 44, 16, 31, -7, 29, -82, 24, 44, 25, 2, 2, 25, -17, 32, 9, -26, -19, -25, 17, -27, 9, -60, 3, 62, -40, -24, -29, -12, 57, 10, -11, 11, -29, -6, 31, -39, 7, -86, 36, 42, 45, 22, -45, 59, -48, 26, 44, 18, -39, -40, 15, -17, -1, -25, -32, 76, -57, -13, -24, -34, 51, 3, 43, 6, -30, -17, -11, -18, -33, -13, 14, 3, -37, -28, -62, 27, -27, -40, 7, 48, 13, -24, -31, -3, -29, -10, 2, 68, -1, -12, -21, -31, 17, 12, 8, 9, 17, -14, -20, -2, 6, -19, 1, 7, 60, -13, -2, 41, 21, -16, -4, 14, -48, -13, -3, 16, 8, -22, -27, 50, -12, -23, -19, -30, 57, -5, 36, 32, -13, -53, -28, 25, -33, 5, 12, 20, 45, -57, -28, 45, -2, -18, 22, -17, -31, 0, -45, 19, 16, -3, 1, -17, -4, -35, 26, -15, 25, -26, 15, 16, -68, -39, -19, 56, -32, 57, -26, 43, 33, -61, -22, 31, 21, -33, -3, -30, -17, 18, 9),
    (53, -7, 49, -17, -20, -3, 9, 17, 23, 21, 44, -6, -33, 13, 8, 16, -2, 28, -6, 22, 32, 55, -38, 34, 28, -1, 23, -3, -1, 49, 0, 22, 52, 16, 31, -13, 3, 6, -6, -6, 8, -28, 11, 15, 0, 7, -13, 1, -15, 4, -26, 35, 49, 68, -3, -12, 17, -6, 46, 1, -15, 12, -6, 16, 7, 13, 9, -75, -25, 6, 4, -3, 20, -6, 23, 1, 28, 8, -19, -12, -15, 1, -24, -15, -26, -3, 35, -6, 22, -41, -22, -23, -16, -28, 6, -20, -18, -69, -19, 27, -20, -22, 15, -18, -11, 56, -29, 11, -43, -49, -2, 6, -4, -5, 25, 16, -13, -12, 16, 8, -25, -4, -3, 16, 26, 23, -5, -45, 38, -55, 5, 41, 18, -6, -29, 9, -27, 47, 52, 14, -70, -1, 20, 67, 25, 32, -12, 26, 28, 33, 16, -22, -27, -28, 1, -16, 25, -14, -3, -27, 31, -46, 31, 21, 18, 26, -37, 49, 19, 21, 49, -19, -67, 11, 18, 42, -15, 60, -26, 13, 5, 41, -21, 9, -24, -18, 5, 20, 2, -5, 21, -12, -21, 0, 2, -41, 4, -7, 5, -34, -3, -65, 39, -19, 34, -11, 12, -32, -20, -16, 11, -35, -9, 34, 39, -35, 23, 10, 14, -24, 20, 25, -26, -35, 4, 51, -49, -92, -26, 11, 33, -17, 0, -75, 23, -36, -12, 0, 46, -13, 22, -46, 46, -42, -14, 27, 21, -6, -5, 18, 12, 20, 28, -31, -23, -25, -49, 3, -25, -31, -4, -1, -3, -36, -69, -46, -7, -26, 2, -13, 23, -19, 9, -90, 50, -36, 10, 14, -9, -16, -36, 40, -16, 22, 49, -30, -48, -4, -6),
    (13, -10, -14, 54, -3, -45, 63, 42, 36, 18, 2, 19, 17, 26, 35, 43, -30, 10, 61, 10, -2, -8, -31, -16, 47, 17, 12, 7, 5, 12, 8, 9, -16, 40, -16, 12, 25, -59, 19, 20, 7, 34, 23, 20, -45, 14, 0, 16, -12, 19, 17, 54, 9, 37, 12, -4, -15, -10, 44, 31, 26, -34, 14, -1, 13, 33, 10, -10, -19, -45, 1, -20, -6, 1, 38, -40, -59, 4, 1, -29, -10, -13, -13, 8, -14, 30, 41, -7, -23, 11, 0, 14, 24, -20, -56, 26, 4, 34, 16, 29, -6, -2, 16, -5, 5, -26, 14, 30, -20, -43, -27, 5, 2, -18, 45, -4, 13, 3, 0, -8, 24, 19, -34, 30, 18, -17, -27, 20, 16, -43, -10, 87, -89, -24, -53, 4, -57, -39, 21, -10, 0, 5, -56, -17, -17, 35, -3, 12, 21, -7, -29, -4, -35, -21, -2, 4, -29, 50, 11, -9, 36, 19, 28, -26, -38, -17, -61, 16, 13, -35, 0, 41, -20, -2, -9, -23, 14, 40, 10, 24, -15, 2, -16, -8, 27, -33, 12, -37, 5, -1, -21, -1, 9, 28, -12, 16, -6, -21, 20, -6, 18, 2, -19, 3, -39, -25, -39, 17, -40, 3, 17, -15, -8, 38, 18, 25, -7, 3, 16, 26, -2, 2, -10, -17, 22, -25, 17, 31, -54, -9, 22, -28, -38, -87, -27, 42, -8, -33, 9, -19, 28, 36, -1, -3, 10, -29, 10, 18, -23, -8, 3, 39, -68, 14, 6, 20, 51, 1, 27, -3, -36, 11, -35, -35, 6, -54, -3, -3, 8, -5, -34, -7, 9, 57, -13, -5, -32, 9, 7, 17, 6, -7, -15, 3, -58, 32, 5, -23, 1),
    (1, -38, -16, 37, -14, 3, 28, -10, 24, -3, 52, 26, -42, -17, 4, -29, 39, 12, -26, -23, 47, 23, 20, 1, 6, -11, 13, 9, 10, 53, 16, -18, -12, -6, 21, 45, -25, 1, -56, -17, -52, -45, 54, 4, -57, -20, -23, -1, 13, -3, -64, -23, 40, 34, 12, 12, 25, -23, 32, -14, -7, 9, -8, -48, -85, 46, -18, 9, 9, -53, -28, 20, -57, 3, 35, -25, -47, 17, -17, 6, -36, -23, -18, 33, 5, 19, 21, -17, 36, 30, -25, -73, 17, -42, 7, 1, 51, 0, -31, 27, -34, 21, 11, -21, 21, -27, 55, 48, -34, -23, -22, -13, 12, -14, -34, -19, 34, 30, 9, 36, -19, -3, 39, -12, 30, 68, 16, -14, 60, -37, 15, 25, -47, 53, -47, 8, -35, -36, 48, 50, -67, -20, -51, -10, 31, 11, -54, -59, 39, -1, 7, 39, -45, 5, 13, 6, 15, 77, -11, -15, 16, -38, -10, 4, -46, 17, -54, 5, -57, -2, 43, 18, -45, 10, -42, 42, -8, 37, -43, -20, 37, 16, 5, -11, -28, 26, -12, 0, 30, 27, -11, -24, -3, 20, -3, 0, -20, -7, -1, -1, 2, -4, 15, 32, -12, -2, -3, -2, -5, -31, -3, 6, -28, 21, -4, 19, 1, -29, 29, 12, -7, 33, 2, 41, 28, -21, -20, -9, -49, 34, -15, 6, -25, -16, -39, 31, -29, 0, 14, 21, 22, -10, -7, -57, 9, -3, -3, 25, -18, 0, -15, 18, -17, 28, -21, 29, 15, -9, -6, 3, -40, 42, -1, 7, -58, -34, -6, 29, -45, -10, -45, -9, -29, 12, 2, -29, 12, -25, 2, -21, -45, 42, 25, 4, -33, 33, -17, 25, -7),
    (-23, -5, -26, -24, 14, 57, 12, 27, -3, 3, -10, -3, -3, -30, 18, -22, 33, -70, 32, -9, -14, -38, 37, 15, -18, -58, 37, 40, 22, 34, 1, -20, -18, -31, -55, 21, 33, 44, 42, 10, 1, -11, 19, -5, 15, -44, 44, -56, 16, -39, -13, 10, -3, -1, 40, 50, -7, -50, 51, 34, 32, -1, -46, -21, -9, 10, -17, -3, 26, -8, -28, -8, -9, -6, 12, 23, -26, 2, 30, -33, 41, 15, -6, -14, -15, -13, -5, 2, -23, 3, 39, 6, 5, -32, -9, -24, -20, 17, -13, 32, 18, 43, 27, 26, -8, 0, -8, 9, 0, 13, 66, -25, -12, -42, 22, 20, -6, -50, 11, 49, -23, 4, 79, -18, -52, -1, -50, -18, -6, 7, -49, -19, 6, 35, 40, 33, -11, 9, 3, 10, 26, 10, 71, -41, 4, -66, -7, 42, 6, 3, 32, 39, -16, -15, -1, 9, -4, 5, -44, -19, -38, 14, -28, -22, -20, 12, -7, 13, -20, -22, -7, -25, 15, -8, 43, -15, 9, -16, 12, 30, 25, 14, 13, 2, -58, -10, 20, 11, -16, 8, -60, -22, 9, 23, -13, 16, 23, -14, 13, 0, 36, 19, -10, 25, 1, 9, 19, -30, 2, -11, -9, 35, -9, -1, -19, -23, -48, 1, 40, -9, 16, -67, -9, -2, -4, 49, -31, -9, 23, 6, -14, 62, 55, 29, 46, -12, 2, -13, 66, -18, 31, -35, -72, 66, 10, 12, 32, -21, -8, -4, 25, 12, 42, -30, 19, 2, -9, 3, -39, -14, 15, -1, -7, 40, 25, 26, 6, -11, 22, -13, 30, -5, -8, -9, -62, 66, 26, 13, 9, -8, -2, -6, -18, 1, 47, 15, -10, -6, 12),
    (-32, 33, -14, 4, 6, -53, 31, 4, 24, 18, 6, -35, 23, 25, 1, 48, -40, 37, 26, 7, -10, 22, -49, -33, 16, 47, 2, -19, -14, -25, 6, 25, 0, 51, 39, -14, 9, -68, 7, 26, 14, -16, 48, -10, 54, 51, 13, 6, -31, 29, 35, 32, 8, 24, -75, -29, 11, 41, -30, -44, -30, -59, 29, -7, 36, 38, 30, 13, 20, -29, -4, -4, 48, 7, 72, -23, 51, 26, 13, -50, 14, 36, -13, 31, 8, 18, 19, -28, -10, 13, -27, -22, -23, -51, -7, -4, -43, 25, -2, 40, 40, -57, 1, 22, 18, -15, -4, 1, 51, 49, 31, 22, -11, -7, 78, 18, -16, 24, -6, -43, -10, 23, -31, -28, -13, -43, -22, -25, -20, 43, 12, 28, 7, -68, 20, 10, 58, 10, 14, -28, 59, 32, 19, 45, -45, 18, 78, 49, -25, 29, -31, 1, -35, 59, -8, -12, -58, -69, 5, -1, -4, 33, -4, 42, -2, -54, -34, -12, 17, 5, 11, -15, 35, -24, 29, 9, -21, -2, 50, 25, -7, 10, -3, -46, -4, -28, -24, -8, 5, -56, 18, -26, 31, 39, 3, 18, 62, -3, -25, -7, 26, 16, 19, -9, 65, 4, 16, 1, -13, -5, 88, 21, -30, -27, 3, -24, -8, 0, 14, -8, -5, -41, -3, -12, -22, 60, 14, -13, 36, -32, 22, 1, -4, 6, -5, 7, 20, 4, 35, 32, -5, 6, 75, -22, 10, -3, -1, 0, -12, 41, -11, -41, -17, -60, 6, 14, -3, 46, -44, -19, -11, 0, -20, 7, 20, -10, 14, 15, 21, -30, 0, -34, -11, 2, 39, 3, -14, -12, 11, 20, -38, 7, 35, -16, 49, -58, 1, 14, -3),
    (30, -42, -24, -13, 48, -9, 38, 10, -1, 43, 12, -7, -30, -28, -4, 50, 11, -32, -30, 11, -3, 29, 27, -23, -20, 46, -38, 14, 44, 12, 7, 9, 21, -67, -41, -25, 23, 37, 32, 8, -13, 20, -47, 19, -36, -71, -44, 25, 2, -52, -18, -12, -35, 10, 41, 39, -5, 43, -74, 42, -15, 35, 37, -1, -6, -40, 22, -2, 6, 32, -6, 33, -9, 15, -18, 24, 9, -20, -21, 14, -7, -40, -3, -39, 23, -5, 21, 4, 0, 18, -3, 42, -3, 55, 10, -5, 22, -69, -30, 2, 3, -39, 0, 14, 20, 15, 12, 3, -28, -40, -29, 20, -32, 11, -7, 27, 0, 71, -12, -40, -49, 24, -13, 20, 7, -13, -12, 8, 41, -30, -7, -37, 17, 6, 49, -10, 43, 41, 5, -9, -44, -59, -10, -10, 28, -6, -8, 6, -5, -3, 72, -6, 0, 28, -56, 66, 25, -18, 22, 5, 33, -21, -4, -30, 16, 17, 12, 10, -15, 11, -27, 9, -28, -79, -3, -21, 5, -18, 14, -54, 8, 16, 67, 1, 24, 9, -27, 58, -1, 6, 5, -10, -2, 8, 1, -11, 23, 6, -26, 22, 7, 7, 41, -3, 11, -3, -14, 11, 10, 49, -14, -17, -13, 29, -14, -15, -20, 16, 30, -39, -16, 15, -11, 12, 8, 29, -27, -26, 9, -13, 13, -4, 54, 2, 8, -28, -10, -8, -13, 10, 13, 45, 13, 17, -2, 56, 10, -44, -43, -25, -4, 2, 32, -51, 14, -4, 21, -2, -30, -28, -3, 39, 1, 15, 35, 13, -6, 35, 0, -11, 18, -44, 9, -7, 0, -11, -17, 21, 31, 1, -19, 12, -14, 17, -8, -19, 9, -9, -5),
    (27, 5, -10, -2, -61, -12, -54, -20, 6, -25, -9, 39, 13, 35, 25, 10, 1, 26, 40, 12, -5, -18, -18, -27, -7, -43, -27, 68, 2, 19, 5, -15, 35, 77, -2, -60, -25, -12, -67, -5, -14, -57, 22, -15, 45, 30, 9, -31, -7, 63, 35, -35, -16, 12, -27, -21, -44, -37, -52, 7, -14, -38, -31, -3, 19, 35, -40, -32, 4, -27, -49, -8, 31, -61, 59, -34, 12, 23, 38, 18, 3, 16, 9, 9, 9, 19, 19, 15, 7, -23, -16, -12, 12, -26, -45, -5, 12, -20, 1, 63, -46, 0, -51, -11, -22, -73, -35, 3, 78, -5, -1, -53, 19, 55, -11, 27, 10, -62, -8, 21, -6, -54, -58, -3, -22, 31, -38, 37, -5, 41, 19, -5, 4, -7, -69, -45, 8, -62, -11, -1, 109, 19, -3, -32, 20, 70, 45, -37, 13, -26, -49, -46, 0, -19, -77, -40, -32, 13, -25, 15, 15, 47, -8, 25, 25, 2, -35, -28, 17, -38, 46, -7, 40, 31, -30, 10, -6, 35, 33, -25, 7, -20, -63, -32, 46, 1, -42, -36, 10, 18, 32, -1, -15, 15, -36, 17, -8, -5, -11, -11, 39, -16, 10, 34, 57, 5, 22, -63, 35, 28, 24, 37, 9, -50, -3, -23, -4, -29, 6, 20, -12, -33, -25, 40, 12, 31, -12, 15, 19, 10, 7, 11, 6, -8, -33, 4, 38, -17, 44, -31, 7, 42, 15, 26, 15, -11, -38, -3, 1, -16, -43, 14, -59, 24, -11, 36, -4, 22, 5, 8, 11, 23, -2, -30, -10, 10, -3, 4, 4, 6, 12, -15, -6, 46, 9, -3, 16, 53, -32, 15, -3, -5, 22, 26, -12, 1, -8, 47, 10),
    (24, -11, 23, 2, 5, -13, -16, 21, 11, 22, 36, 22, -51, -11, 27, -33, -12, -2, -16, -14, -21, 5, 28, -16, -22, 0, 43, 2, 13, -38, -11, 7, 48, -18, 11, -12, -4, -20, -24, 15, -31, 39, -38, 29, -71, -31, -50, -39, 25, 7, -44, 15, -43, -6, 25, 13, -8, -5, 15, 23, -7, 5, -7, 11, 34, -21, -6, 19, -25, -2, -34, -3, -49, 2, -15, 1, -5, -3, -52, 20, -16, 16, -48, 14, -8, 21, -39, -24, -8, -5, 21, 16, -14, -5, 14, 2, 56, -34, 29, 13, 20, 1, 50, 35, 12, 57, 46, 63, -78, -25, -33, -29, 24, -17, -79, -40, 17, -5, 43, -3, -12, 12, -11, 52, 61, -21, -3, 20, 69, -79, 31, -59, -5, 73, -12, 15, -24, 66, -32, 43, -56, -33, -65, 46, 29, -15, -44, -38, 30, 32, 63, -6, 7, 25, -55, 63, 14, -21, -8, -6, 28, -20, 2, -26, -12, 35, -53, 11, -37, 20, -18, 34, 20, 10, -11, 21, -2, 23, -23, -18, -15, 53, -3, -10, 25, -17, -50, 43, -30, -12, 7, -14, 24, -2, -8, 1, 1, -14, -5, -2, -4, 13, 20, 34, -19, 3, -41, -3, 7, 13, -39, -37, 14, 12, 27, -23, 27, 10, -11, 26, 29, -12, -21, 48, -1, -36, 0, -53, -8, 15, -37, 1, -40, -6, 6, -22, -17, -4, -13, 33, -26, 0, -20, -26, 19, 54, 34, -32, 21, 42, -29, 9, 9, -42, 22, -3, 3, -22, -4, -33, -8, 13, -10, -20, -19, -3, -52, -38, 7, 13, 29, 50, -19, 5, 17, 20, -18, 24, -20, 3, 6, 4, 4, 16, 3, -13, 22, -14, -2),
    (-15, -10, 13, -19, 28, 5, -6, 50, -7, -4, -37, 20, 68, 18, 24, 39, -49, -7, 29, 53, 6, 35, -7, -27, -3, -5, -8, -5, -43, 14, -34, 18, 12, 7, -1, -37, 8, 8, 31, -1, 7, -11, -48, 20, 65, 42, 56, 57, -52, -1, 25, 42, -37, 44, -11, -13, 19, -35, 35, 13, -54, -35, -24, 33, 9, 26, -23, -28, -20, -22, 5, -22, -27, -30, -27, 0, 14, 21, -21, 15, -54, -3, 28, -14, -9, 32, -1, -38, 26, 15, 10, -6, -17, -15, 2, 34, -24, 36, 37, 1, 26, -32, 7, 41, 31, -1, -31, -26, 54, -4, 0, 29, -35, -10, 23, 47, 3, -8, -39, 18, 16, 8, -23, -33, -7, -5, 4, 16, -45, 36, 15, 18, -7, -46, 41, 63, 18, 52, 10, -35, 38, 36, 5, 98, -23, 26, 0, 73, -9, 29, -42, 2, 18, -23, 63, -25, -55, -34, 3, -3, 40, 32, 54, 9, -30, -62, 21, 24, -7, 51, 20, 20, 16, 38, -24, 62, -31, 36, -29, 49, -8, 34, -29, -19, -4, -6, 4, -12, -19, -20, -12, 15, -27, 10, 13, -8, -2, -30, -10, -37, -13, 0, -31, -2, 18, -22, -10, -33, 24, 16, 19, 0, 9, -41, 21, -23, 3, 10, -8, -41, 14, 22, -12, 0, -32, -1, -21, -13, 13, -46, -19, -4, 1, 22, -21, -28, -40, -17, 25, 1, 4, -1, -7, 10, 5, -17, 11, -8, -21, 2, 4, 15, 39, 25, -10, -1, 15, -3, -12, 10, -1, -42, 21, 45, 21, 43, 15, -3, -25, 5, 18, 38, -21, 13, -26, -2, 8, -25, 27, -21, -24, -31, 9, 16, 49, -17, -9, 33, -8),
    (20, -17, -38, -48, 9, -5, -23, 21, 26, -37, 43, 33, 44, 4, 18, -28, -18, -27, 23, -38, -18, 22, -8, 21, -48, -30, -67, -7, 20, -67, -4, 33, 25, 47, -33, -18, 39, -25, -3, -8, 72, -22, 76, 9, 43, 41, -39, 30, -61, -38, 61, 17, 10, 2, -17, 0, -18, 0, -78, -39, 31, -49, 3, 9, 20, 65, 27, -19, 20, -66, 20, -13, 24, -10, -7, -9, -55, 36, -9, 18, -3, 15, 27, 0, -10, 2, -10, -20, 20, 8, -14, -9, 14, -38, 35, 12, 12, 62, 16, -66, 39, -44, -13, 11, 43, -17, 53, -14, 45, 12, 17, -17, -34, -14, 38, 4, -5, 14, -2, -22, -30, 25, -44, -20, 52, -78, 2, 44, -5, 98, 20, -73, 41, -82, 13, -7, 67, 27, 50, -25, -13, -3, -53, -9, -32, 11, 67, -28, -8, -23, -3, -10, 11, 23, -20, -3, 41, -62, 48, 21, -42, 49, -18, -10, 2, -35, 30, -16, 34, 22, 17, 14, -25, -45, -21, 12, 3, -12, -12, -49, -40, 6, -19, 7, -6, 35, -12, 27, -16, -4, 50, 20, 9, 32, -12, -34, 12, -9, 12, -8, 25, 20, -13, 7, 19, 38, 4, -4, -3, 3, 26, -38, 12, -13, -27, -11, 17, -21, 12, -5, -7, -2, -6, 64, -1, 44, 4, -2, 21, -45, 51, 21, 17, 34, 18, 7, -40, 6, 2, -12, -20, 1, 49, -36, -28, -8, -43, -11, 11, 7, -12, 4, 21, -17, 26, 45, -7, -7, -32, 37, 0, 32, 9, -1, 8, 17, -24, 17, 34, -58, 8, -38, 6, 0, -63, 42, -13, 1, 4, -40, -17, -8, -6, -10, 21, 34, -12, 0, -8),
    (-29, 8, 14, 34, -30, 7, -9, 2, 31, -22, 4, -21, 44, -21, -17, -13, 7, -2, 3, -7, -22, -11, -9, -29, 3, 26, 46, -2, -22, 16, -11, 3, 1, -17, -4, 0, -35, -25, -38, -1, 34, -35, 39, -47, 16, 23, -8, -22, -2, 12, -8, -3, 27, 18, -11, 22, 13, 11, 12, -88, -7, -19, -31, 27, -15, 26, 4, 26, 10, -26, 11, 10, 14, -6, 63, -40, -30, 21, 2, -29, 0, 32, 0, 35, 54, -3, -9, 15, 5, -4, -4, -45, 48, 2, 23, 31, 10, 51, -11, 29, -21, -6, -72, -31, -16, -18, -17, -14, 66, -23, 20, -20, -28, 27, -19, 7, -37, -38, -49, 12, 14, -35, 24, -64, -33, -22, -13, -10, 8, 40, -3, 30, -2, -68, -35, -3, 25, -2, 74, -32, -1, 96, -18, 14, 15, 40, -4, 21, 35, -16, -74, 18, -19, -19, 7, -85, -8, -6, 3, 84, -2, 68, -27, 29, 38, -43, 20, 22, 28, 9, 74, 26, -71, 38, -16, -30, 19, 5, -2, 8, 18, -23, -18, -28, 19, 4, -8, -37, 46, 22, 5, 31, 24, 2, -4, 11, -22, 0, -28, -11, -19, -18, -25, -24, 7, -5, 5, -5, 34, 24, -30, 21, -16, -1, -46, -17, -33, -85, 61, -9, -49, -14, -1, 4, 33, 10, 8, -5, 8, -41, -14, -5, -15, 12, 10, 18, -8, 53, -24, 33, -1, 53, -11, 5, -12, 18, -86, 30, 11, -37, 31, -6, -15, -4, 4, 62, -23, 22, 9, 1, 10, -11, 2, 10, -18, 14, 34, 24, -40, 16, -8, -18, 1, 29, 22, -13, -27, -12, -18, -17, -22, -23, 36, 7, 27, -1, 14, 20, 1),
    (-2, -6, -4, -4, -53, 48, -3, 6, -35, 13, -28, 1, 18, 11, 34, -1, -15, -1, 1, -44, 23, -24, -6, 47, -30, -6, -54, 3, -12, -4, -61, -15, -13, -10, -9, -21, -31, 74, -16, -43, -28, -23, -21, 11, 15, 11, 30, -41, -16, -4, -4, -18, 14, -25, -26, 41, 2, 27, -4, -10, 2, -17, -62, -26, -14, 26, -19, -9, -43, 84, -6, -57, 22, -3, -22, -17, 14, 30, 39, -19, 12, -6, 26, 21, 8, -6, -55, 3, -9, -2, 15, -32, -31, -28, 0, -6, -5, 11, -27, 28, 17, 30, 9, 27, 2, -3, 89, 11, -29, 11, 27, 23, 40, 10, -19, -4, -26, 40, 30, -20, -50, -23, -23, 14, 80, -18, -29, 16, 22, 12, -25, 11, -11, 48, 4, 17, -6, 9, 97, -21, -12, 0, 33, -10, 23, 13, -4, -26, -12, 24, 31, 19, 13, 4, 19, 9, 88, -13, 7, -14, -27, 4, 9, 28, 11, 11, -2, -31, -5, 7, 26, 5, 37, 1, -41, 10, -19, -18, -1, 13, 48, 32, 31, -43, -27, 26, 30, -18, 28, -13, -5, -19, 5, -16, -42, 6, -14, -2, -31, -11, -1, -41, 18, -15, 18, -6, -4, -15, -17, -5, -2, 7, 14, -20, -40, -36, 30, 34, 31, -48, -5, -10, -31, -3, 32, 14, -46, -7, -14, -4, -21, 7, 11, -22, 64, -29, 23, -11, -6, 7, 14, -7, -44, 2, 40, -11, -26, -7, 21, 32, 26, -55, 52, 10, -6, 14, -10, 32, -7, 26, 2, -22, -24, -5, 6, -4, 22, 4, 0, 4, -25, -6, -19, -25, -51, 14, 46, 22, 5, -1, -9, 53, -47, -31, 28, 5, -28, 12, 14),
    (22, 2, -20, -16, -33, -25, -110, -17, -16, -35, 15, 0, 41, 62, -29, -15, 1, 64, -44, 34, 10, -20, -41, -11, 12, -4, 2, -15, -25, -19, -59, -8, 10, 46, -4, 18, -21, -39, -47, 8, 34, -28, 56, -24, -32, 55, 37, 12, -35, 58, -15, 24, 0, 36, -15, -23, -10, -3, 10, -20, 21, -44, -5, 39, -20, 40, 17, 7, 2, -22, -14, 27, 44, 15, 5, -6, -18, 34, 40, 21, -35, 43, -25, 2, -9, 34, 0, -6, 14, 14, 4, -12, 0, -4, 21, 38, 18, 19, 16, 40, -14, -26, -40, -9, -15, -33, -2, 10, 8, 33, 3, 5, 0, 84, -34, 9, 4, -46, -38, -16, 25, -72, 49, 6, -81, 1, -18, 74, 36, 72, 23, -25, 22, -11, -14, -30, 18, -3, 48, 25, -37, 42, -71, 27, 9, 84, -5, -43, -17, 21, -17, 26, 6, -32, 58, -9, -2, -15, 20, 78, 34, 37, 33, -10, 3, 11, 18, -17, -3, -13, 18, 31, -57, 17, 10, 49, -13, 29, -2, -10, -26, 51, -44, 6, -19, 0, 62, 11, -23, -50, 1, 30, 27, -1, 13, 1, 24, -12, -8, 18, 10, -23, 7, -1, 20, -47, 18, 1, 25, 42, 15, 16, -21, 25, 13, 8, -20, -27, 33, 5, -25, -2, 6, 48, 12, -9, -10, -39, 5, 33, -15, -30, -11, -26, -19, 36, 29, -40, -27, -41, 20, 21, -46, -30, -3, -7, 25, 6, -4, -17, -23, -6, 23, -17, -6, 11, 15, 1, -15, -54, 6, 24, 4, -45, -24, -16, -2, 32, -58, -33, 4, -98, -16, -7, -28, -30, -11, -8, -10, 7, -45, 28, 0, -11, -29, -48, 14, 19, -4),
    (-25, 9, -51, 35, -4, 18, 28, -30, 6, -32, -59, 1, 27, -16, 2, -36, 25, -7, 13, -50, 7, -36, -3, -30, 17, 4, -10, -2, 6, 7, -24, 23, -17, -3, -18, -49, 15, 26, 35, -6, -5, -10, -79, 0, 13, 29, -18, -23, -17, -38, -1, 16, -7, -27, 22, 4, 51, -38, 20, -9, -3, 18, -31, 27, -36, 15, 14, -47, -35, -3, 12, -6, -16, -2, -53, 29, -5, 18, -38, 28, -50, -74, -21, 21, -61, -27, 19, 23, -2, -43, 8, -6, 23, 22, -4, 29, 7, -3, 25, -22, -8, 42, -27, -9, -4, -39, 1, 12, 26, 40, -62, 17, -33, 1, -30, 14, 74, 5, -6, -8, 19, 6, 43, -58, -21, 10, 4, 19, -26, 15, 35, -20, 10, 13, -1, 4, 9, -18, -50, -32, 33, 69, -44, 36, -29, 3, -52, 93, 68, 31, 13, 16, 27, 26, 24, -40, -67, -13, -18, 39, -8, 11, 35, -11, 2, -25, 7, -10, 33, -27, -19, 6, 36, 40, 34, 1, -15, 1, -40, 57, 0, -36, -2, 24, -24, -5, -35, -2, -22, -26, -5, 43, -9, 31, 27, -6, -43, -2, -25, 24, -33, -6, -14, -21, -18, 8, -39, -11, -35, -14, -32, 9, -16, -35, -10, 1, -37, 52, -6, -37, -34, -21, 18, -21, -29, 40, 3, 10, -12, -44, -16, -11, 16, 4, 23, -40, 2, 3, -6, 32, -24, 49, -29, 64, -9, 1, -16, -36, -2, 47, 37, -64, -4, -47, 34, -19, 32, 38, -3, 6, -3, -21, 17, -14, 27, 11, 10, -6, -11, 37, 39, 27, -7, 29, -60, 60, -17, -13, -22, -10, -23, 44, -22, -22, -8, -51, 31, -26, 1),
    (-30, 79, 45, -96, 35, -8, 3, 25, 14, 14, 32, -23, 31, 26, 32, 28, -13, 5, 23, -5, 19, 8, 13, -22, 16, 4, -79, 2, 15, -40, 0, 4, 10, 41, 1, -77, 52, 24, 35, 17, 84, 34, 2, -27, 27, 73, 43, 9, -6, 23, 21, -5, -38, -11, -15, 13, 20, -21, -65, -20, 39, -44, 1, 17, 17, 13, -24, -33, 32, 24, 17, -6, 56, 40, 1, 28, -49, 29, 31, 13, -22, 13, -3, 50, -37, 5, 0, -17, -32, 7, 13, -2, -18, -25, -2, 30, 33, 45, 5, -78, 18, -23, 19, 31, 14, 17, 17, -13, -19, 42, 0, -6, -5, 6, 46, -39, 14, -3, -67, 10, 15, 10, -21, -16, 15, -19, 41, 21, 6, 35, -5, -58, 15, -54, 34, 7, 61, -20, 36, -19, -39, 4, -8, -24, 10, -21, 38, -42, -37, -4, -23, -36, 7, 33, -53, 38, 36, -42, 21, 38, 0, -26, -1, 23, -48, -13, -21, -9, 50, 3, -18, 8, -52, -25, -15, -7, 31, -22, -3, -23, 70, -39, 3, -25, -9, 0, 4, 0, -8, 44, 6, -14, -41, -43, -10, -21, -11, -39, 53, 2, 35, -1, 19, 7, -37, 28, -38, 3, -33, 24, 20, -22, -32, 5, -35, -7, 34, 11, -7, -15, -11, 24, 19, 27, -36, 4, -3, 9, 8, -18, 21, -29, 18, -3, -15, 2, -25, -28, 23, -8, -4, -29, -24, -23, 15, -12, 34, -38, 33, 51, 15, -28, 3, 46, -21, 33, 12, -54, -11, 5, -28, 25, 46, -6, -2, -7, -26, 14, 6, -7, -41, -5, 6, -24, -4, 0, 6, -36, 6, -18, -30, 28, 12, 16, 6, 24, 1, 17, 0),
    (-13, 24, 6, -37, 12, -17, 37, 21, 21, 5, 4, 32, -33, -43, -40, -5, -44, -46, -20, 15, 21, -35, 45, -17, -15, 8, 36, 24, 38, 21, 28, 21, 11, -16, 23, -14, -6, -5, -17, 14, 2, 18, -17, 38, -55, -50, -48, 4, -35, -6, -46, 14, 4, -28, 45, 20, 17, 13, 14, 21, 31, 46, 15, 5, 1, -9, -13, 18, 16, -1, -37, 11, -20, -25, 3, 8, -28, -6, -3, -32, -7, -6, -24, -19, 4, -37, -17, 29, 2, 3, 1, 20, 19, 28, 25, 20, -16, 9, -17, -25, 18, 10, 37, 39, 28, 42, 14, 12, -58, -46, -10, 27, 8, -37, -29, -4, 23, 46, 69, 11, 21, 58, 56, 20, 40, 6, -15, 4, 3, -51, 21, -15, 20, 12, 19, -1, 36, -1, -18, 53, -53, -42, -33, -10, 14, -19, -11, -22, 2, 1, 94, -3, 29, -22, 8, 59, -12, 10, -21, -6, 35, -55, 41, 49, 10, 5, -46, 18, -8, -41, -73, 55, -19, -3, -37, -29, 19, 2, 4, -8, -3, -38, -4, -18, 0, -59, 6, 20, -12, 25, -29, 19, 43, -21, -2, -14, 8, -27, 6, -10, 8, -6, -1, -14, -21, -37, 13, -34, -37, -7, -42, -4, -3, 4, 34, 19, -32, 22, -33, 1, 11, -6, 7, 3, 20, -37, 26, -48, 7, 17, -10, 24, 39, 18, 2, 35, -35, -32, -37, -1, -17, -32, 29, 5, -7, -4, 37, 26, 20, -3, -25, 3, 30, 3, -46, 27, 26, 1, 7, 10, -1, 8, -12, 36, -21, -1, -29, 6, 29, 17, -36, 7, 19, 21, 7, 27, -18, 7, 13, -21, -9, -66, 1, 1, 17, -17, -41, 18, -5),
    (3, -5, -17, 4, 2, -36, -11, 10, 0, -7, -29, 0, 1, 16, -9, -19, -10, 21, -45, 19, 52, -23, -49, -28, 41, 1, 14, 19, -8, -25, 24, -1, 9, 57, 31, -48, 7, -41, 22, 56, 0, 17, 38, -6, -54, 19, 3, -17, 13, 3, -58, -35, 17, 44, -19, 8, 41, -34, 48, 18, 40, -8, -3, 62, -17, 11, 6, -15, 15, -22, 0, 26, -16, 24, 53, -12, -24, -23, -18, 15, 22, -69, 5, -35, -31, 17, 14, 46, 8, -3, 42, 53, 5, 21, 1, 60, -19, -1, 10, -8, 9, -15, -47, -38, -27, -19, 30, -32, 23, 4, -11, -34, -11, 26, -71, -6, 38, 3, 12, 3, -63, 57, 52, -70, -19, 6, -18, -42, -28, 40, -12, 24, 6, 10, -60, -26, 21, -43, -8, -45, -1, 29, 4, -35, 8, 21, -37, 7, 8, -38, -11, -58, 11, 20, -16, -70, 25, -23, -17, -26, 11, 5, 24, -35, -27, -28, -32, -1, 8, 8, 8, -38, -18, 71, 11, -5, -35, 14, -11, 12, -28, -9, -33, -29, 17, 33, 6, -31, 36, -19, -24, -1, 22, 15, -16, -1, -32, -11, 31, 25, 3, 18, 25, 13, 13, 35, -23, 35, 8, -17, -10, 10, 1, -12, 29, 25, 17, 10, -45, 6, 3, 3, -4, 18, 28, 17, 3, -54, -14, -4, 10, -21, -31, 4, 31, 1, 26, -5, -19, 42, -12, -3, 6, 11, 1, 18, 5, -6, -21, 10, -33, 35, 25, -12, 27, 17, -13, -17, 12, -54, -5, 17, -9, -34, -9, 0, 19, -36, 44, 2, -17, -14, 1, 49, -37, -42, 35, 31, 21, 16, 12, -8, -61, -15, 2, 8, 18, -10, 3),
    (46, -8, -13, -60, -6, 22, 30, 15, 15, -21, 23, -12, -31, -22, 16, -28, 49, 32, -18, -43, 1, -4, 17, -15, 8, -40, 8, 64, 32, -7, 24, 20, 53, 23, -29, -3, 6, 3, -13, -40, 12, 5, -12, 19, 5, -53, 3, -38, -7, 38, 14, -13, -24, -21, 24, -43, 1, -61, -11, 48, -31, -23, -6, 3, 27, 6, -20, -15, -26, 2, -38, -40, -41, 13, -24, 15, -19, -28, 67, 11, 21, 12, 38, 18, -23, 8, -9, -5, 12, -29, -15, 46, -23, -27, 4, 15, -6, 5, -52, -3, 16, 93, -44, -8, -16, -26, 20, -1, 39, -47, 14, -34, 2, 1, -14, 8, 18, 18, 17, -27, 15, -35, -24, 9, -19, 10, -10, -15, -17, -31, -32, -36, 11, 25, -28, -8, -3, -1, 6, -33, 92, -9, 39, 14, 20, 12, -11, 24, 0, 54, 1, -32, -30, -42, -68, 6, -28, -20, 50, -5, -3, -20, -43, -38, 16, -4, 34, -12, 2, 4, -6, -39, 25, -19, 46, 14, 8, 3, 8, 51, -33, 22, 7, -19, -7, -4, -21, 40, -5, 1, 33, 0, 5, -18, -31, 1, -5, 36, -32, -3, -9, -11, 17, -15, 67, 33, 41, 38, 26, 53, 5, 41, -36, 29, -10, -38, 6, -3, 16, 6, 14, -71, -30, -53, 8, -23, 15, 8, -3, -28, -10, -12, 18, 22, 22, -2, 57, 48, 13, 39, 1, 31, -30, 35, -9, 5, -71, -35, -6, -4, -20, -52, 3, -7, 30, -10, -30, 18, -6, 9, 33, -12, -2, 1, 8, 36, -16, -34, 36, 44, 15, 41, -12, 39, -1, 30, -6, 29, -21, -2, 36, 9, 1, -31, 11, -6, 32, -25, -6),
    (-1, -35, 18, 32, 3, 27, 3, -11, -22, -18, 46, 18, 26, -29, -23, -32, -49, 16, -9, 23, 27, 7, -29, -5, -40, 27, -27, -63, -24, 31, -5, -10, -12, -8, 20, -18, -4, 16, -13, -11, 18, -2, 2, -2, 32, 34, -31, -26, -4, 8, -17, 4, 48, -11, -1, -6, 6, 56, -28, -82, 31, 33, 17, -1, -4, -16, 40, -17, 7, 13, -8, 23, 32, -1, 35, -18, 31, 46, -7, -10, -4, 18, 7, 23, 20, 11, 0, 33, -12, 15, 3, -53, 30, 29, -4, -20, -44, 28, -7, 34, -37, -24, -15, 2, 21, 9, 49, -6, -14, -28, -17, 1, 19, 40, -31, 1, -20, -8, 0, -9, -48, 20, 7, -1, 46, -12, 21, 24, -14, 45, -23, 40, -5, 37, -14, -15, 34, -19, 10, 3, 83, -5, -67, 8, -44, 47, -21, 20, 31, -65, -74, -10, -46, 52, -13, -109, 25, 44, -32, -13, -14, 57, 9, 17, -3, 14, 4, -6, 21, -4, -15, -38, 28, 22, -25, -19, 15, 45, 13, 21, 51, -48, -61, -11, -17, -10, 6, -46, 43, 49, -12, 0, -24, 63, 8, 28, 8, -27, 8, 15, -12, -26, -1, -21, -14, -47, -9, -6, 9, 2, 5, -19, -34, -27, -29, -3, -7, -28, 20, 6, 50, -6, 5, 1, 10, 21, 19, 32, -47, 31, 19, -9, -45, 6, -45, 5, 10, -4, -58, -36, -49, 20, -23, 32, 4, -71, -84, 3, -10, 20, 45, -45, -58, 33, -26, -16, 8, 45, 25, 53, 5, 4, 13, -7, 26, 17, -26, 18, 62, 5, 11, -12, -24, 23, -3, -8, -15, -46, -60, -2, -9, 8, 26, -32, -12, 18, 36, 19, 6),
    (-23, -58, 5, 22, 13, 9, 31, 3, -14, 60, 44, -13, 14, 23, -10, 52, 28, 51, -34, 21, 19, 55, -5, 33, 24, 28, -26, 15, 7, -8, 10, -39, -8, -27, 13, 46, -6, -3, -16, 8, -56, 24, -8, 4, -24, 18, -62, 16, 0, 6, -47, -10, 56, 6, -24, 55, 24, 23, 39, -23, -11, 13, -7, -19, 38, -29, 30, 34, -36, 1, -13, 11, -22, -8, 0, -15, -16, 7, 23, 36, 6, 37, -50, 5, 55, -25, 10, -1, 3, 28, -7, -39, 13, 28, 9, -7, 2, -33, 32, 9, -53, 26, -5, 40, 3, 7, 24, -7, -37, 23, -37, 25, 17, -1, -16, -25, 16, 15, 13, 23, 23, 23, 8, -10, 31, 8, -17, -52, -19, -38, -3, -17, -47, -32, -20, -6, -29, -21, -9, -30, 3, 25, -50, 31, 7, -27, -42, -16, 24, 24, 0, 38, 3, 38, -33, -55, -21, -26, -14, -28, -12, 38, 22, -54, -25, -39, -5, -9, -28, -19, -35, 12, -1, 18, -17, -30, 9, -20, -48, -26, 12, -29, -14, 21, 6, 5, 6, -29, -6, 13, -1, 39, -24, 5, 29, -5, -5, -3, -13, -45, -18, -18, -2, -18, 3, 6, -72, -6, -29, -8, -10, -46, 28, -2, -12, -7, -7, 13, 7, -11, -1, -19, -36, -9, 1, 46, 31, -22, -14, -21, -17, 16, 4, -20, 4, -24, 9, 43, -43, 3, -28, -48, -35, -20, 36, -23, 28, 3, -29, 40, -43, -82, -34, 17, 14, 25, 14, 7, -11, -3, 7, -41, 25, 15, 8, 0, -33, 6, -9, 11, -36, -4, -27, -31, -26, -22, 12, 29, -12, 31, 6, 6, -2, -59, -6, -19, 46, 7, -6),
    (47, -30, 21, -42, 28, 8, -6, -2, -24, 16, 46, -10, 15, -13, -7, 2, -60, -45, 17, 33, 29, -5, 1, 2, -13, 18, -2, -26, 13, -34, -49, 35, 22, -1, 23, -32, 11, -61, 42, -8, 9, -7, 32, 19, -30, 13, -26, 24, -27, -2, -4, 12, 12, 18, -50, -8, -3, -15, 19, -17, 26, -27, 30, 58, -4, 13, 31, 12, -2, -27, 9, 5, -16, -39, 28, -5, -58, -16, -69, 0, -19, 37, -35, -24, -4, -4, -4, 4, -12, 3, 22, -3, 2, -8, 16, 53, 6, -2, 14, -16, 3, -59, 19, -5, 25, 11, 33, 59, -57, -22, -87, 15, -64, -41, -39, 6, 17, -11, 52, 31, 27, 28, -6, 5, -6, 6, -7, 43, 39, 61, 20, 3, -15, -70, 34, -10, 52, 6, -4, 81, -69, -57, -70, -6, -9, -63, -33, -40, -29, -36, 44, 3, -19, 35, -23, 65, -27, 11, 16, 72, 13, 14, -10, -29, -33, -15, 28, -7, 13, -15, 2, 51, 12, -37, -2, -4, -8, -51, 23, -70, -28, 3, 1, 22, -18, 42, 27, 3, 11, -11, -15, 69, 19, 25, 29, -23, 23, -11, 28, -6, -13, 32, 29, 47, -29, -52, -2, -25, -9, -14, -15, -7, -11, 22, 50, 16, 38, -5, -48, 24, 11, 22, -11, 60, 19, 43, -27, -26, 8, 18, 18, -5, 47, 4, -34, 26, -16, -15, -58, -10, -5, -33, -18, 8, 18, 1, -6, 16, -13, 24, 0, 15, 0, -9, -26, 31, -14, 7, -28, 1, -10, 8, -5, -6, 14, -23, -7, 29, -21, -1, 2, -3, -10, -41, -22, -9, 13, 6, 11, 0, 41, 45, 0, -60, 2, -56, -11, 31, -7),
    (-20, -3, 3, -16, 8, -12, 26, 23, -2, -8, 1, 13, 15, -4, 17, 39, -32, -19, 28, 0, -14, 28, -7, 18, -16, 26, -15, 16, 8, -26, -34, -11, 6, -39, -33, 2, 9, 2, 37, 7, -20, 24, 37, 1, -23, -9, 46, -2, 26, -23, 20, -28, 15, 28, 43, 30, -1, -2, -7, 21, 27, 33, -22, -27, 13, -34, -6, 8, -10, -1, 1, 8, -36, 6, -26, 31, -12, -36, 34, -22, 28, -45, -12, -64, 8, 15, 16, 17, -7, 0, 10, 29, -4, 56, 11, -15, -43, 16, -18, -25, 44, -18, 19, 28, 32, 39, 64, 13, -44, -1, 42, 2, -9, -51, -17, -20, 19, 56, 19, -29, 12, 65, -53, -22, 33, -24, -35, 29, -6, -39, -40, -41, 17, 29, 14, 15, -31, 29, 22, 19, -37, -53, 6, -12, -17, -75, -6, -61, 30, 10, 68, 22, -21, 31, -30, 13, 39, 49, -31, 2, 9, -47, 14, -22, -3, 40, 21, -2, -1, 14, -8, 42, -32, -23, -18, -28, 14, -44, 31, -47, 14, -41, 46, 16, -14, 5, -28, 35, 10, 34, 13, 3, 19, -20, -65, -4, 38, 11, -1, 15, 22, 0, 33, 14, -50, -37, 31, -19, -22, -43, -19, -49, 12, 19, 26, -34, -19, 23, 13, -36, 59, 3, -52, 19, 13, -31, -36, -23, -7, 50, 25, 10, 7, -11, 16, 60, -34, -39, -4, -61, 5, -39, -15, -17, 41, -29, 33, -21, 28, -16, -38, 38, 0, 52, -21, 9, 41, -12, 13, -36, -7, 26, -5, -5, 20, -4, -16, 32, -17, -7, -7, -36, 9, -23, 21, 21, 5, -22, 26, 3, -1, -8, -17, 18, 17, 16, -13, 30, -4),
    (-34, -41, -2, 54, -22, -16, -9, -30, 27, -19, 48, -21, -73, -68, -17, -14, 21, -21, -12, -21, 18, 18, 65, -14, 0, 31, 21, 10, 51, -5, 12, -59, -41, -21, 17, 22, 1, -20, -22, -4, -46, 6, 26, -41, -23, -49, -3, -23, 33, 17, 8, -12, 9, 21, 52, -42, -8, -5, 21, -6, 35, 0, -5, -21, -12, -11, 10, 40, 3, 11, -37, -33, -36, -14, -10, -10, 12, -17, -14, -16, 21, -22, 45, 17, 2, -15, -2, -6, -6, -26, 24, -43, -6, -32, -10, 5, 12, 14, -21, 28, -24, 13, -20, 8, 21, -7, 52, 25, -51, -37, 17, -60, -14, -33, -48, -33, 28, -26, 27, -12, 18, 26, 44, -14, 30, 20, -38, 11, 19, -6, -32, 63, -40, 14, -23, 20, -18, 26, 39, -3, -57, -45, -26, -30, 12, -49, -76, -57, 65, -39, 69, 4, 26, -24, 24, 17, 63, 56, -26, 16, 14, -18, -2, 24, -9, 12, -62, 18, -36, -4, 17, -10, -10, -50, -7, -13, 8, -61, -57, -7, 52, -25, 21, 24, -12, -8, 0, 7, 38, 34, 3, 24, 16, 25, -7, 18, -10, 27, -37, -2, 6, -36, 4, 32, 16, 14, 24, -16, 5, 9, -14, -9, 3, -15, -17, -7, 3, 8, -10, -45, 4, 19, -7, -5, 33, 19, -7, -20, -14, 39, -14, 27, -18, -27, 4, 36, -12, 9, 24, -37, 22, -7, 2, 28, 19, -45, -13, -7, -8, -15, 11, -36, 59, 68, -30, 7, 21, 7, 14, -16, -2, 17, -25, 28, -23, -22, -39, 14, -13, 17, 17, 1, -18, -11, -17, 4, 22, -15, -4, 17, -42, 7, 10, -27, 18, 39, -15, 19, 1),
    (31, -46, 6, 38, -16, 29, 18, -4, -51, 47, 10, 41, -96, 9, -2, 10, 38, -3, -8, -45, -23, 26, -17, 42, 12, 11, -32, 54, -7, 19, -12, 0, 24, -23, 13, -3, -49, 44, 18, 29, -58, 23, 23, 38, -103, -35, 5, 34, 47, 3, -41, -70, -10, 62, 12, 25, -13, -3, 13, 73, -7, -11, -1, 9, -9, -15, 37, 2, -38, 26, -15, 22, -22, 9, 20, 11, -53, -41, -19, 21, 1, -12, -36, -71, 22, 44, 18, 24, 2, 7, 1, 11, -7, -4, -16, 16, 35, -24, -15, 5, -36, 21, 17, -8, -59, 0, 1, 20, -34, -43, 41, -30, 38, -25, 25, -94, -15, -15, 21, 20, -24, 4, 5, 44, 14, -9, -44, -13, 27, -12, -23, -53, -35, 50, 15, -23, -64, -31, 4, 16, -52, -30, 35, -40, -4, -17, -1, -102, -18, 4, 34, 54, -44, 7, -7, 41, 37, -17, -30, -31, 16, -1, -13, -49, -18, 29, -11, -4, -25, -71, -15, 10, -38, -19, 18, -25, 19, -15, 2, -89, -11, -4, 4, 24, -25, 9, 22, 33, 11, -25, -17, 1, 1, 12, -22, -54, 29, 4, -13, -23, -3, -8, -44, 13, 27, -6, 42, 5, 23, 6, 28, -15, -51, 19, 2, 3, -16, -4, 36, -22, 16, 19, -52, 8, 5, 6, -11, -44, 1, 6, -7, -12, 33, -48, -49, -16, 25, 19, 85, -12, 39, -11, 29, -34, -22, -5, 29, 1, 7, 10, -17, 12, -10, -11, -23, 6, 30, 15, -3, -41, -25, -1, 21, -12, 8, -40, -6, 1, -31, -6, 34, -12, 23, -17, 3, -37, -14, -35, 47, 1, 31, -54, 5, -13, -22, -11, -21, 26, -11),
    (-38, 10, -43, 43, -8, -7, 4, -39, -18, -46, -14, -10, 19, 17, 3, 12, 12, -18, -72, -18, -16, -19, -24, -13, -10, -45, 24, -41, 24, 28, -33, 31, -25, 32, 16, 74, -11, -45, -5, 26, 5, -35, -25, -18, -17, 27, 5, -2, -29, 43, -35, 26, -27, -9, -4, -37, -2, -43, 50, -33, 8, 31, -23, 32, 8, 11, 4, 44, -24, -23, -23, 27, 2, -32, -15, 26, -9, 7, -17, -18, -4, 29, -24, 0, 11, -9, 13, 10, 13, -16, 50, 5, -26, 28, -7, 47, -29, -17, 15, 56, 5, 4, -13, 53, -46, -2, -27, -20, -35, 17, 0, -9, 35, 30, -32, -5, -11, 15, -30, 22, 26, -68, 60, -18, -29, 2, 33, 19, -15, -27, 50, 62, -2, 8, -21, 51, -41, 27, 31, 10, -28, 3, 29, 10, 31, 63, -31, -5, 40, 31, -5, 41, 42, -42, 32, -23, -44, 18, 4, 8, 9, 4, 39, -7, 14, 28, -16, 36, -33, 1, 49, 5, 6, -3, -15, 16, 30, 29, -19, -2, 60, 8, 19, 8, -6, -8, 13, -12, -34, -5, -9, 2, -18, -15, -14, -15, 7, 12, -14, -17, -16, 6, 43, -30, 27, -27, -2, -26, 22, -20, -39, 23, -7, 22, 61, 0, -32, 17, 13, -14, 24, -22, -26, -19, -30, -34, -35, 24, 15, 9, -2, 2, -55, 2, 27, -60, 13, -20, 5, -24, -6, -10, -21, 7, 20, 19, 42, -10, -23, -2, 7, -27, 39, 15, 2, -52, -7, -11, -45, 32, -1, -9, -9, -46, -18, 8, 41, -49, -19, -20, -7, -18, -13, -8, -27, 4, 24, 1, -44, 8, -41, 13, 16, -19, -7, 30, -6, -32, -4),
    (-16, 13, -24, -17, 10, -12, 10, -24, -8, 27, -11, 10, 45, -21, -26, -14, -9, -7, -21, -25, -6, -68, 17, -1, 12, 16, 35, -33, 37, 5, -42, 30, -31, 12, 11, 64, 26, -28, -16, 0, 4, 31, 10, 8, 30, 2, -29, -22, -55, -41, -11, 50, -7, -32, -11, 30, 9, 19, 1, -29, 21, -13, -14, -7, -10, 5, 15, 9, -2, -16, 6, -7, -23, 11, 34, -33, 24, -29, 20, -10, -20, -30, 22, 37, 27, -17, -6, 24, 6, -28, 53, 9, -1, -2, -9, -2, -43, 17, -24, 24, -31, -11, -6, -18, 2, -59, -59, -29, 30, 22, -42, 13, -12, -23, -65, 32, 29, -13, -11, 15, -13, -19, 29, -26, -24, 2, -25, 15, -9, 26, -43, 40, -14, -55, -1, -37, 1, -28, -13, -37, 37, 24, -25, 24, -46, -11, -67, 52, 41, 20, 6, -23, 26, -3, -4, -35, -10, 26, -18, 16, -37, -13, 15, 31, -18, -47, -22, -9, 32, -37, 30, -28, 38, -14, -2, -23, -17, -36, -24, -6, 22, -9, 38, 8, 25, -36, 7, -37, -2, 64, -23, 29, 1, -7, 14, 99, -19, 8, 21, 1, -27, 22, -44, -9, -6, 24, -30, 37, 3, 45, -13, 59, 0, -17, -30, 8, 13, -50, -15, -15, -56, 53, 30, -15, 2, -23, 17, 74, -22, 11, 4, 53, -9, 15, -12, -9, 4, -2, -5, 30, -8, 48, -40, 52, 0, 15, -57, -7, 12, -61, 78, -30, -37, 13, 57, -16, 17, -6, -10, -10, 10, 8, -4, 43, 28, -34, 0, -2, 38, -16, 6, 3, 13, -22, -39, 22, 11, 29, -29, 14, 11, -41, 5, -4, -8, 20, -14, -11, -1),
    (3, 10, 24, 7, -16, -73, 19, -13, -9, -6, -18, 27, -15, 4, 7, -18, 34, 55, -51, -17, -37, -3, 6, -7, -3, -62, 26, 10, 1, -25, -14, -3, 43, 50, 7, 40, -33, 9, -30, -2, -23, 6, -7, 37, -41, 20, 41, 40, 7, 55, -62, -26, -11, -33, 7, -8, -2, -25, 54, 10, -6, -5, -8, 22, 3, -1, -2, 39, -36, 50, -27, -8, -22, 11, 18, 35, -25, 49, -8, 0, -13, -4, -53, -39, 15, -22, -1, 32, 37, -1, -11, -30, -18, -24, 18, 1, 17, 35, 30, -28, -3, 6, -57, 18, -27, -8, -12, -6, -11, 36, -43, -6, 0, 32, -37, -25, 5, 18, -3, 6, 25, 22, 10, -1, -3, -2, -5, -13, 30, 15, 45, -82, -41, -21, -76, -23, -64, -64, -28, -16, -78, 52, -27, 39, 24, 29, -60, -32, 15, 39, -6, 27, 46, 13, 4, 0, -20, -45, -24, 27, 36, 23, -8, -23, -33, -14, -25, -27, -51, -28, -18, -32, -11, 43, 21, 43, -18, 26, -31, -29, -12, 30, 5, 11, 18, -4, 21, -4, -33, -21, -10, 31, 41, 30, -12, -52, 9, 22, -17, -25, -18, -64, -23, 38, -14, 21, -31, -3, -3, 2, 19, -14, -10, 10, 7, -17, 9, 8, -11, -7, -16, 5, 14, 9, 73, 4, 21, -43, -32, 24, -40, -46, -16, -50, 1, 27, -38, 32, -32, -1, 35, 8, -13, -44, 29, 42, -28, 4, -5, 13, 0, 5, -33, 28, -7, 18, 65, 22, 47, -34, -5, 5, -40, -14, -14, -47, 0, 41, -21, 36, 18, 1, 0, 35, -6, -43, -12, 15, -39, -1, 6, -23, 56, 7, -10, 15, -28, 31, -1),
    (20, -16, -21, 66, 16, -31, 26, -39, 18, -21, 29, 2, 5, 41, -22, -11, -13, 28, 8, 11, -32, -6, -47, 8, -26, -69, 40, 17, -38, -35, 11, 47, -15, 32, -22, 23, 27, 7, 28, 10, 32, 31, 10, 13, -28, 29, 8, -13, -12, 18, -29, 13, -35, -12, -31, 19, -17, -42, 31, 1, -4, -30, 7, 65, -64, 20, -42, 9, 55, 0, 7, 15, 37, 0, 49, 15, -11, -2, 16, -8, -28, -24, -27, 10, -65, -14, 4, 6, -12, -14, 53, -8, 40, -27, 5, 47, -46, -46, -4, 98, -2, -52, 7, -20, -3, 9, 33, -2, 50, 13, 10, -5, 19, 27, 37, 58, -19, 20, 3, -50, 38, -43, 43, 3, -25, 7, 12, -43, 37, 18, -35, 66, 7, -49, 36, -13, 12, 16, 29, -1, 38, 35, 81, 28, -2, 17, 36, 17, -34, 33, -6, 2, -14, -66, 30, 20, -70, -18, 48, -9, 22, 52, -17, 17, 12, -29, 37, -18, 37, 1, 10, 12, 37, 26, 50, -6, -31, -9, 19, -1, -41, -27, -39, 18, 5, -28, 17, 35, -6, -63, -1, 48, -11, -22, 9, 14, -15, -3, -46, 25, 36, 12, 31, -11, 39, -31, -111, -30, -2, -32, -27, -40, 41, -12, 24, -29, 13, 4, -13, 0, 61, 52, -26, 5, -15, -34, 3, 74, -12, -10, -7, 0, -10, 30, 30, -38, -2, -31, -22, -27, 3, -23, -35, 10, 47, 5, 16, -19, 4, -8, -5, 17, 17, 69, -19, 5, -41, -4, 6, 46, 0, -34, 12, -37, 14, 7, 10, -20, -28, 29, 17, -19, -31, 23, -4, 17, -48, -19, -7, -24, 1, -41, 24, 13, -38, 42, 55, 12, 3),
    (14, -35, 14, -13, -25, 20, -37, 27, 7, 16, -29, 33, -91, -21, -13, -42, 10, -2, -6, -39, 16, -14, 15, -13, -18, 12, 25, -10, 33, 1, 42, -8, 26, -44, 58, -11, -15, 39, -30, 46, -30, 28, 23, 11, -95, -13, -11, 33, 5, 9, -47, -12, 47, 32, 47, -18, -9, 4, -12, 0, 19, -23, -3, 14, 24, -1, 25, -12, -2, 47, -19, 34, -11, 13, 24, 43, -37, 20, -44, 36, 20, -15, -40, -32, 41, 52, 33, 5, -22, 4, -5, 15, -14, -38, 12, 11, 3, 10, -24, -13, -2, -11, 12, -30, -13, -34, 13, 18, 0, -7, 15, -40, -11, -50, 19, -57, 7, -31, 2, 4, -11, 41, -26, 31, 23, 8, -38, -27, 22, -45, -46, -70, -37, 34, -22, -52, -32, -26, 3, -2, 16, -28, 23, -11, 14, -68, 4, -39, -11, -29, 34, 31, -3, 62, -62, 20, 8, -7, -42, -69, -32, -17, -3, -50, -40, 45, -17, -46, -25, -19, -10, -41, 13, -5, 14, 10, 10, -82, -16, 12, 13, -5, 24, 18, -53, 12, -23, 9, 26, -18, -28, -52, -10, 73, 4, 6, 14, -26, -21, -20, -23, 11, 37, -43, -22, 29, -29, -6, -22, 17, -9, 12, 8, 43, 1, 17, -3, 52, 3, -7, 36, -17, -16, 41, -21, 34, 35, -4, 8, -3, -37, -9, 23, -3, 18, -10, -37, 16, -38, -36, 9, 7, 3, 5, 0, 39, 37, -18, -12, 25, 26, -27, 22, 20, -30, 25, -1, -3, -6, -12, -1, 3, -14, -42, 20, -33, 19, -12, -22, -2, -1, -24, 10, 24, -24, 13, -1, 13, -18, -56, -9, -14, 30, -25, -17, 1, -45, 13, -1)
  );
  ----------------
  CONSTANT Flatten_1_Columns : NATURAL := 4;
  CONSTANT Flatten_1_Rows    : NATURAL := 4;
  CONSTANT Flatten_1_Values  : NATURAL := 48;
  ----------------
  CONSTANT NN_Layer_1_Activation : Activation_T := relu;
  CONSTANT NN_Layer_1_Inputs     : NATURAL := 768;
  CONSTANT NN_Layer_1_Outputs    : NATURAL := 10;
  CONSTANT NN_Layer_1_Out_Offset : INTEGER := 3;
  CONSTANT NN_Layer_1_Offset     : INTEGER := 0;
  CONSTANT NN_Layer_1 : CNN_Weights_T(0 to NN_Layer_1_Outputs-1, 0 to NN_Layer_1_Inputs) :=
  (
    (-11, -23, -6, 0, 3, -27, -9, -21, -15, 1, 13, 2, 11, -12, -20, -15, -15, 3, 19, -27, -15, -7, 26, -11, -17, 3, -1, -12, -20, 0, 18, 7, 14, -19, -13, -3, -20, 29, 4, -4, -10, 24, -11, -7, 14, -12, 2, 4, -28, 8, 6, -11, -3, -34, -9, 21, -14, 6, 6, -3, 20, -11, -2, -25, -7, -6, -1, -33, -25, 10, 36, -19, -37, -5, -6, -4, -15, -8, 10, -27, 16, -1, -2, 1, 1, 6, 2, -3, -22, 23, -30, 10, 11, -21, 35, -8, 5, 12, 2, -13, 18, -17, -1, 16, -15, 6, 0, 11, 20, -5, 33, 13, 3, 0, 4, 10, 2, 6, 14, -11, -7, -7, -7, 14, -16, -9, 3, -25, -2, -12, -2, -4, 27, -2, 15, -18, -18, 11, -9, 9, 8, -10, 25, -4, 14, 10, -14, -13, 14, -16, -15, 12, 10, 14, -10, 4, -9, 4, -1, 21, 4, 5, 11, -3, 0, 7, 11, 5, 4, -3, -12, -15, -5, -1, -8, -5, 23, -4, -9, 1, 3, -21, 8, -12, 8, 3, -32, 5, 7, 14, 4, -15, -13, -25, -21, -13, 0, -21, -12, 5, -25, 25, 3, -9, 39, 10, 4, -12, -27, 1, -9, 4, -12, -34, 12, 12, -29, 12, -27, 0, 18, 14, 21, -4, 21, -11, -30, -5, -19, 21, -13, 5, -40, 29, -20, -8, 13, -10, 37, -30, 4, -37, 0, -21, -23, -36, 4, 60, -29, 21, 9, -15, 35, 9, 10, -27, -42, 4, -33, 16, -17, -12, 28, -25, -44, 2, -26, 5, 12, 9, 17, -11, 19, 0, -31, -3, 10, 26, -22, 8, -50, 37, -26, 0, -2, -22, 65, 2, 6, -31, 1, -11, -20, -14, -1, 45, -36, 6, 26, 1, 15, 6, -9, 2, 11, -2, -37, 6, -20, 12, 36, -70, -41, 8, -21, 6, -9, 4, 10, -16, 6, 3, -2, -1, 18, -23, 1, -2, -42, 21, -22, 0, -4, -10, 49, -21, 5, 0, -8, 4, -6, -7, -18, 13, -20, 18, 1, -15, 0, 4, -3, 10, -8, 0, -5, -3, -7, 20, 15, -11, -10, 8, 19, -18, -16, 0, 21, -3, -2, -3, 2, -6, 11, -1, 14, 8, -27, 16, 6, 4, -9, 5, 23, -20, -5, -21, -9, -32, 2, -15, 2, 21, -19, 1, -4, 7, 0, 9, -2, -1, -7, 6, -7, 4, -4, -56, -5, 8, -27, 9, -13, 2, 16, 11, -1, 10, 20, -14, -20, 5, 15, 7, -13, -8, -44, 3, -4, 5, 11, -10, 19, -2, 6, -60, 3, -37, -1, -28, 11, 22, -34, 8, -3, 22, 21, 20, -1, -8, -5, 23, -32, 2, 15, -17, 11, 15, -40, 4, -12, 12, 18, 18, -7, -4, 7, -5, -20, 6, 8, 0, -21, 8, -61, 30, -9, -5, 21, -2, 32, 6, 2, -64, 3, -22, -8, -9, 2, 34, -30, 0, 13, 36, 17, 11, -15, 6, 23, 6, -51, 8, 6, -8, 20, 7, -60, 4, -2, 7, 1, 2, 15, -8, -6, 6, -1, 6, 8, -14, 0, -18, -12, 17, -10, 14, -4, -17, 31, -8, 11, -19, -42, 13, -14, -7, -17, 17, 0, 14, 6, 12, -5, 2, -7, 5, 6, 8, -14, -5, -3, 4, 23, -4, -34, -9, -19, -3, 18, 12, 21, -17, 0, 7, 0, -24, 14, -26, 2, -48, 1, 4, 31, 20, 5, -3, -6, 7, 1, 5, -9, -10, 12, 10, 1, 7, -11, -7, 0, -2, 10, 4, -8, 10, -9, -6, -4, -2, -10, 10, 9, -13, -10, -16, -7, 1, 3, 6, 2, 3, 3, -11, 4, -2, -1, -1, -3, 3, -7, 17, -7, 4, -7, -3, 6, -16, 12, -33, 6, -37, 6, -27, -2, 10, -13, -4, -4, 12, -11, 2, 1, 6, 17, -4, -21, -8, -7, 7, -5, -9, -16, -8, 8, 12, -5, -6, -4, 6, -15, -16, -9, 9, 8, -13, -22, -19, -9, 18, 0, -10, 8, 9, 5, -2, -9, -5, 0, -11, -3, -35, 5, 6, -8, -16, 8, 15, -3, -17, 8, 0, 15, 13, -13, 4, 8, -8, 17, 0, -27, -10, 5, 0, 13, 5, 8, -9, 10, 4, -2, 3, -2, -3, 2, -30, 8, 11, 3, -5, -2, -13, 12, -12, -1, -1, -55, 6, -6, 1, 0, -8, -14, -23, 10, 9, 13, 12, -6, -2, -3, 5, 0, 8, -3, -2, 2, 7, -8, -11, -16, 10, 10, 3, 13, -6, -9, 2, -24, -16, 5, -17, -10, -17, -3, -1, 4, 8, 6, 2, -17, 6, 4),
    (-11, 21, -11, 16, 11, -9, -5, 1, -6, -20, 3, 12, -44, -9, -27, 27, 26, 9, -22, -31, 12, 8, 16, 11, -1, 7, -34, -38, -10, -11, 14, -5, -18, -11, 11, -32, 10, -3, -28, -17, 13, 10, -17, -20, 1, -20, -2, -19, -49, 33, -15, -7, 14, -6, 0, 0, -28, -18, 3, 5, -31, 10, -31, 18, 14, 9, -9, -20, 39, -13, 25, 26, 8, 11, -14, -16, 11, -45, 18, -27, -1, -7, -6, -31, 1, -5, -36, -34, 10, -2, -55, -36, -2, -38, -10, -11, -38, 19, -14, -2, 5, -19, -4, 3, -27, -21, 4, 2, -19, -5, -1, 4, 13, 5, 18, -5, -2, -25, 5, 10, 6, 23, -12, 10, 8, -11, 9, 5, -5, -8, -18, -15, 0, 5, -25, -12, -1, -13, -35, -21, -8, -15, 19, -4, -1, 9, -18, -12, -10, -22, 6, 5, -5, -7, 12, 5, -1, -14, 4, -11, 10, 1, 2, 2, 0, -30, 3, 11, 10, 2, -18, -21, 12, 7, 7, 6, -2, -6, -9, 5, -3, 15, -9, -12, -13, -26, -13, 0, 0, -1, -9, 4, -21, 36, 1, 11, 9, 4, 11, 6, -22, -10, 32, 5, -21, 25, -13, 33, 39, 9, 11, -36, 16, 3, 17, 25, 8, 18, -36, -39, -13, -17, 7, -46, -19, -9, 18, -25, -5, -3, -21, -53, 3, -4, -21, -10, -14, -27, -8, -11, -42, 56, -11, -13, 18, -16, 21, 1, -46, -29, 32, -7, -37, 62, -27, 16, 29, 23, 30, -22, 40, -12, 55, 45, 7, 23, -20, -12, -3, -62, 9, -58, -17, 6, -15, -31, 8, 2, -6, -72, 15, 28, -62, -26, -15, -22, -16, -57, -31, 34, 3, -13, 2, -9, 23, 0, -15, -28, 34, -10, -21, 9, 1, 16, 25, 11, 32, -7, 13, -15, 25, 25, 8, 36, -7, 4, 14, -34, 5, -25, 2, -4, -30, -16, 9, -8, -4, -40, 25, 2, -22, -32, -11, -7, -2, 1, -24, -7, -24, -8, -3, -6, 0, 1, 3, -24, 3, 3, -5, -5, 3, 10, 7, -13, 1, -2, 9, -31, 4, 6, -5, -1, -15, -6, 23, -6, -15, -22, -11, 1, -9, -1, 10, -7, -9, -4, 4, -12, -5, -2, 1, 1, -5, 18, -17, 21, 0, 13, 9, 2, 21, -6, -16, -15, 18, 4, 1, 12, -12, 19, 16, 8, 5, -2, 3, -1, 8, -15, 5, -1, 9, -25, 12, -19, -4, -42, -7, 1, 1, -32, 2, 1, -37, -19, 18, 12, -11, -15, 4, -26, 5, -9, -42, 34, -21, 0, 12, -18, 14, 12, -15, -18, 21, -13, -34, 36, -23, -1, 31, -11, 24, -4, 19, 1, 17, 5, 14, 6, 6, -13, 0, -43, 2, -48, -17, -5, -14, -31, -4, -11, -18, -39, 28, 2, -44, -24, 7, -31, 9, -20, -21, 19, -11, 2, 1, 1, 3, -8, 7, -29, 26, -1, -12, -10, -11, 1, 5, -6, 27, -15, 28, -13, -5, 17, 27, 9, 11, 4, 14, -11, 10, -25, -2, -6, -14, -12, -6, 12, -6, 9, 17, 5, -10, -25, -2, -26, 1, -7, -12, 9, -16, -17, -2, -3, -3, 10, -9, -10, 7, 4, 21, -12, -7, -8, 5, -22, 6, -13, 2, -15, 6, 9, -1, -5, -8, -19, 15, 17, 7, -16, 4, -1, -6, 0, 4, -8, -28, -33, 8, 0, -45, -16, 7, -32, 0, 6, 5, 20, -9, 12, -6, -5, 11, -5, -14, -1, 9, 2, -27, -9, 2, 7, 4, 7, 6, -3, -6, -11, 11, 1, -4, 1, -13, -20, -7, -11, 9, -28, -10, 5, -5, -4, 2, -1, -9, -9, -4, 1, -16, -8, -1, -15, -5, -1, -21, 16, -14, 12, 8, -10, 10, 4, -15, -2, 0, -3, -26, 6, -12, 13, 4, -10, 9, -15, 4, -2, 2, 5, 6, -6, -7, -12, 0, -11, 2, -30, -20, -5, 3, -17, -2, 11, -5, -18, -1, -7, -20, -10, 3, -29, -20, -8, -11, 12, -17, 7, -6, -25, 6, -5, -14, -1, -5, 12, -12, -6, 2, 9, -10, -9, 12, -16, -2, -19, 1, 10, 4, -14, -11, -8, -6, -15, 7, -29, -6, -10, -1, -20, 12, 6, -15, -3, 12, -1, -13, -3, 2, -26, -2, 9, -11, 6, -46, -23, 2, -22, 6, 11, -29, 3, 12, -2, -8, -14, -5, 6, 7, 0, -1, 0, 9, -6, 12, -5, 0, 9, -12, -21, 4, -19, -6, -15, -2, 5, 8, 13, 4, -7, -7, -25, -7, 4, 9, -13, 12, -20, -3, -5, 6),
    (-39, 12, 14, 12, -12, 12, 11, 12, -10, 17, -2, -20, -1, -9, -25, -2, -10, 9, -28, -12, -11, -1, -13, -10, 9, -8, 15, -1, -17, -12, -18, -33, -9, -6, 20, -8, -24, -7, 7, 12, 10, -9, -1, 0, -20, 1, -2, -6, -62, 11, 14, 3, -7, 24, 5, 11, -1, 17, -18, -18, -1, -9, -22, 5, 12, 27, -39, -13, -29, 5, -13, -25, -10, -16, 3, -14, -23, -32, -36, -21, 19, -35, 28, -14, -24, -7, -1, 10, 30, 0, 1, -20, -31, -10, -17, -35, -34, 5, 6, -3, 20, 19, 8, 5, -21, 24, -22, -5, -14, 2, -19, 0, 5, 14, -18, -9, -20, 8, 10, -18, -9, -20, 1, -16, -34, -9, -21, -14, 30, -38, 11, -17, -3, 1, -9, 13, 43, 4, 9, -9, 4, -27, -9, -18, -7, 2, -3, -9, -5, 3, 4, 2, 0, -4, -5, 5, -21, -1, 0, -1, 6, 7, -6, -6, -8, -1, 8, -1, -18, -8, -23, -11, -5, -20, -1, -6, 2, -15, 1, -6, -3, -16, 2, 5, 21, 2, -2, 5, 7, -12, 4, -1, -40, 5, 2, 32, -11, 9, 35, 19, -17, 15, 1, -37, -2, -41, 18, 9, 1, 21, -9, 8, -1, -22, 5, 3, 10, -29, 13, -18, -9, -5, -14, -18, 13, 0, 18, -3, -35, 7, 7, 8, 11, -4, -26, 11, -21, 1, 5, -12, -51, -8, 8, 24, -26, 22, 37, 18, -20, 3, 14, -14, -10, -50, 31, -33, 33, 34, -6, 14, -15, -9, 2, 17, 1, -33, 17, 10, -7, -25, -53, -15, 28, -10, 18, -2, -47, 15, 0, 6, 21, 0, -41, 4, -31, 0, 10, -10, -38, -5, 9, 12, -7, 10, 41, 6, -15, -2, 11, 3, -13, -10, 19, -20, 19, 13, -24, 6, -32, 13, 1, 16, -17, -36, 22, 23, -17, -26, -51, -40, 31, -8, 8, -12, -43, -1, 3, 4, 15, 9, -29, -7, -11, -6, 6, -7, -13, -10, -2, 5, 5, 21, 25, 5, -6, -7, 7, 6, -21, -3, -10, -21, -1, -8, -8, -4, -13, -2, -1, 7, 2, -24, -18, 13, -2, -13, -21, -9, 25, -21, 0, -17, -9, -2, 0, -11, 15, 5, 4, 2, 5, -13, -11, 10, -18, 4, -21, 5, -1, 3, 1, 10, 0, 9, 0, -10, -17, -25, 1, -5, -13, 0, 16, 12, 28, -20, 0, 21, 0, -31, 8, 4, 11, -9, -10, -9, 17, 2, 4, 5, -20, 3, 9, -6, -3, 6, -27, 7, -10, -3, -10, 1, -23, 1, -1, 12, 5, 11, 18, 15, -4, -3, 7, -7, -1, -24, 17, -42, 36, 23, 20, 16, 6, -22, -10, 22, -7, -29, 25, 19, 27, -16, -31, -14, 30, -1, 2, 9, -27, 22, -3, 2, 4, 10, -22, -9, 6, 1, -21, 9, -25, 7, -8, 0, 6, 3, 15, -15, 10, -4, 6, 11, -5, -1, 19, -28, -17, 8, 15, 4, 10, 0, -21, 24, -16, -6, 20, 24, 21, 4, -30, -16, 35, 2, 12, -3, -28, 18, -2, 6, -12, -9, -31, -1, 5, 1, -6, 16, -18, 3, 15, -2, 7, 6, 0, -4, 1, -14, -11, 1, 6, -2, -6, -11, 4, -3, 4, 6, 15, -8, -6, 11, 11, -10, 7, 21, 3, -12, -21, -1, 14, -1, -1, 10, -10, 1, -5, 19, 9, 4, -10, -21, 1, -14, 7, -6, 2, 3, -5, 5, -11, -7, 11, -6, 12, 5, 1, -13, -11, -15, -5, 0, -12, -3, 4, 0, 0, -4, 10, 4, 3, 0, -6, 7, 15, -5, -22, 13, -2, -7, -11, -10, -18, 21, 15, -2, -3, 8, -13, 10, 5, 13, -8, 2, 0, 7, -6, 9, 4, -12, 2, 3, 15, -9, 9, -9, 3, -37, 12, -21, 6, -2, 13, 11, 1, -14, -9, 6, 0, -10, -16, 8, 16, 2, -4, 5, 18, 2, 6, 6, -13, 18, 14, 10, -9, -7, -4, -11, -2, -4, -22, 11, -1, -2, -1, 17, 12, 8, -5, 2, 14, 12, 5, -12, -2, -26, -3, -13, 1, 6, -14, 0, 4, 4, -10, 8, 2, -2, -16, -9, -11, -15, -7, -2, -7, 6, -1, 8, -10, -5, -4, 19, -5, 9, -8, -7, -13, -2, -9, 6, -10, 6, 35, -5, -1, -8, -1, 1, -4, 2, -8, 3, -1, -9, -8, -5, -11, -6, 5, 8, 2, -2, -12, 8, -3, -16, 12, 8, 5, -9, -10, -22, 1, -8, 2, -1, 2, 4, -5, 19, 12, 2, -6, -13, 8, -5, -5, -6, -3),
    (2, -15, 24, -16, -18, 15, 18, -4, -2, 23, -2, -21, 5, 12, -13, -6, -14, -14, -22, -16, 14, 22, -7, -3, 14, -36, 14, -17, -41, -26, -13, -21, -3, 3, 25, -1, -1, -16, 8, 16, 15, -2, 27, -12, 5, 0, 1, -4, 16, -19, 5, -15, -20, 32, 2, 3, 10, 10, -7, -16, 9, 17, -11, -6, -4, 12, -28, -16, 5, 19, -10, -15, 21, -8, 5, -14, -44, -45, -13, 2, -5, -29, 34, 8, -3, -32, 15, 5, 28, 9, 30, -11, -11, 10, -8, -11, 22, -3, 3, -17, -16, 24, -13, -10, 9, 12, -12, -11, -8, 15, -5, -1, -19, 3, -21, -22, 2, 6, -5, -18, -4, -9, 14, -29, -31, -32, -10, 6, -2, -24, 28, 0, -19, -12, -1, 2, 9, 12, 26, 0, 3, 12, -6, -2, 5, -1, 7, -4, -15, 0, 1, -8, 3, -7, 4, -7, -6, 4, -2, -6, -8, 17, -15, -14, -1, 16, -5, -13, 8, 2, 3, -25, -7, -8, -3, 13, 1, -5, 2, -8, -9, 4, 10, 1, -13, 12, 2, 6, -8, 1, 4, -2, -3, -21, 29, -17, 20, 7, 2, -19, 11, 13, -5, -24, -9, 15, -14, 0, 16, -10, -59, -18, 19, 29, -15, -4, 13, -19, 13, -11, -25, -18, 4, -4, -22, -6, 25, -9, -3, -30, 12, 6, 15, -9, 17, -15, -14, 1, -6, -11, 11, -36, 14, -7, 24, 23, -17, -16, 7, 2, 5, -40, 4, 15, -19, 14, 23, 1, -51, -22, 24, 26, -34, -19, 30, -9, 6, -9, -37, -31, -15, 2, -29, -18, 11, -7, -3, -35, 14, 4, 24, 3, -2, -16, -13, 11, 6, -38, 20, -24, 17, -9, -1, 15, -33, -10, 19, 1, -13, -22, -2, 14, -37, -2, -6, 0, -31, -18, 4, 15, -23, -17, 19, 6, 6, -16, -42, -25, -15, -2, -43, -9, -1, -7, -8, -20, 6, 6, -1, 1, -2, -17, -5, 9, -4, -21, 18, -6, 0, 8, -14, -6, -8, -8, 2, 2, -3, -21, -6, 2, -15, -3, 6, -3, -15, -20, -1, 11, -3, -11, -2, 2, 10, -2, -24, -3, -14, 18, -9, -12, 0, -4, -9, -3, 12, 5, -6, -3, 4, -1, -2, 17, 6, -9, -14, -37, 25, -7, 9, 3, -1, 14, -8, 9, 5, -2, 2, 17, -11, -15, 0, -15, -30, 0, 12, -6, 1, 11, 3, -5, 11, -22, 3, 4, -24, -3, -32, 0, 17, 1, -4, -24, -6, 15, 14, -1, 12, -11, -3, -3, 6, -16, 8, -42, 24, 2, -1, 6, 2, 5, 3, 6, -2, -12, 17, 16, -1, 19, 3, -14, -42, -6, 1, 12, -12, 0, 12, -9, 15, -5, -15, -5, -16, 3, -22, -4, 12, 2, 8, -28, 2, 9, 15, 3, 4, -8, -6, 2, -2, -26, 20, -23, 10, -1, -17, 3, -13, -2, 6, 5, -13, -25, 12, 9, -5, 8, -8, -13, -24, -4, -1, 4, -2, -11, 33, -9, 17, -11, -15, -11, -9, -3, -38, 2, 9, 0, 15, -32, 1, 13, 7, 1, -3, -13, -4, -3, 2, -17, 23, -12, 8, 18, -3, -6, -10, -11, 10, 8, -12, -18, 14, 3, -7, -3, -7, -10, -10, 6, 1, 7, 5, -10, 14, -6, 1, 5, 1, 3, -4, 5, -19, 2, 7, 8, 2, -4, 15, 6, -2, -11, 12, 0, -5, 20, 4, -6, -8, -13, 21, 13, -9, 2, -3, -5, 0, 23, -8, -9, 4, -5, 0, -15, -30, -4, -11, 5, 0, -7, -3, -1, 8, -7, 3, -9, 7, -2, -7, 7, -15, -2, 18, -12, -8, -8, -2, 7, 20, -5, 5, -1, -1, 2, 5, 6, 2, -28, 18, 1, -9, 1, -8, -1, -4, 10, -7, -4, 10, 8, 1, -2, -25, 6, -14, -4, 8, 1, -5, 10, 8, -7, 18, 1, 4, -14, -4, -5, -4, 11, 6, -1, -1, -1, -18, -6, 15, -7, 6, 13, 8, 1, 7, -1, -15, -11, 8, -4, -15, 3, -14, -4, 8, -1, -1, -11, 10, 17, -14, -16, -31, 2, -12, 3, 1, 2, 4, -9, 10, 8, 19, -6, 7, -20, -17, -2, 9, 12, 11, -11, 6, -2, 5, -16, 16, -12, 5, 7, -7, 7, -3, -5, 7, -4, -11, 17, -15, 3, -6, -16, -14, -3, 3, 1, -11, -2, 7, 3, -10, -8, -16, -6, -6, -2, -8, 3, 10, -15, -3, -4, -14, -6, -10, -8, -12, -10, -6, 5, 8, -13, -17, -2, 12, -14, 6, -5, 8, -11, -13, -14, -11),
    (17, -7, -8, -37, -5, -25, 6, 18, 21, -26, -15, 20, -39, -6, 45, 4, 1, -10, -19, 50, 2, -3, -6, -2, 1, 1, 12, 21, -4, -12, -18, 25, -10, 5, -15, 3, 28, -28, 5, -10, -28, -36, -15, 9, -2, 8, 3, -8, 15, -9, -20, -48, 34, -13, 9, 12, 22, -61, -19, 27, -29, -16, 51, 8, 0, -18, 16, 37, -5, -4, 18, 14, -2, -8, 0, 25, -30, -16, -13, 24, 17, -41, -31, -8, 14, -17, 5, -33, -29, -28, -19, 28, 9, 12, -5, -25, -14, -6, -29, -13, -18, -21, 12, 11, -17, -52, -16, 26, -8, -11, 23, 1, 20, -6, 1, -1, 3, -17, -6, 5, 0, -5, -12, 31, -30, -14, -18, 9, 20, -22, -36, -4, -1, -13, 9, -44, -8, -27, -13, 4, 1, 13, -7, -9, -20, 1, -28, 3, -7, -14, 5, 5, 8, -3, -13, 14, -4, 0, 6, -15, 1, 0, -5, 8, -10, -12, -12, -5, 12, -10, -35, 3, -3, -9, -15, 0, -1, 10, -6, -1, -7, 0, 13, -29, 7, -17, 2, -15, 17, -8, -3, -1, 17, 3, -7, -25, -8, -9, 1, -1, 19, -39, -30, 54, -13, -12, 24, -24, -24, -15, 19, 30, -4, 5, -2, -30, 21, -13, 21, 24, 15, -23, -24, 5, -5, 4, -13, 1, 32, -30, 11, -11, -2, -51, 28, 7, 14, 19, -11, 43, -3, 17, -12, -39, 11, -9, 0, 3, 21, -44, -43, 60, -12, -16, 36, -4, -29, -17, 18, 32, -10, -2, -2, 8, 28, -13, 16, 18, 1, -26, -17, 8, 1, -10, -2, 12, 29, -29, 9, -10, 4, -49, 30, 21, 29, 17, -19, 68, -14, 17, -10, -16, 11, -1, 6, 1, -4, -38, -33, 44, -11, -4, 17, 0, 0, -14, 4, 15, -7, 13, -17, 30, 15, -16, 8, 7, -15, -18, -18, -10, 15, -8, -3, -1, -4, -20, 14, -36, 18, -33, 26, 3, 9, 13, -27, 36, -16, 10, -5, 9, -8, -12, 11, 4, 6, -14, -9, 31, -18, 8, 10, -3, -9, -4, 13, 0, -3, -1, -5, 7, 6, -7, -48, 17, 9, -13, -15, 2, 24, 2, -17, -16, 1, -17, 6, -15, 14, -19, 10, 6, -6, -4, -17, 0, 3, 29, -24, -13, -6, -16, -34, -17, 33, -12, -22, 6, -1, -5, 11, -14, -3, 3, 22, 7, -11, 24, 8, -13, 18, -13, 14, 19, -7, -32, 23, -5, -10, -14, -8, -2, 5, -5, 20, 16, 1, -21, 23, -2, 4, 10, -20, 33, -7, 35, -30, -17, 7, -17, -31, -17, 42, -21, -39, 18, -4, -29, 12, -27, -9, 0, 20, 0, -36, 0, -21, -16, 15, -3, 8, 11, -17, -24, 7, -5, -13, -19, 10, -2, -15, -19, 18, 8, 9, -23, 36, 8, 9, 19, -40, 42, -20, 33, -16, -8, 5, -2, -12, -24, 29, -24, -24, 6, -16, -18, 14, -5, -18, -15, 9, 2, -15, 7, -28, 2, 30, -8, -12, 1, -11, -5, 0, -7, -6, 0, 4, -24, -9, -5, 23, -3, 11, -4, 24, 5, 13, 15, -30, 37, -6, 0, 8, 0, 13, -8, 7, -12, -1, -14, -4, 0, -11, -1, 13, -13, -12, -1, 8, 5, -7, 8, -8, 13, 10, -3, -2, 14, 12, 1, 3, -9, -8, -3, 0, 7, 0, -9, 0, 5, 3, 2, 12, -5, -8, -24, -9, 14, 5, 0, -19, 11, 1, -1, 6, -3, -2, -14, -2, -5, -12, -6, 16, -7, 10, -4, 15, -2, 2, 16, 4, -2, 3, 12, 21, 0, -7, -8, -10, -14, -28, -9, -5, -6, 0, 4, 16, 5, -4, 4, 24, -5, 3, -2, -1, 13, -6, 5, -36, -11, -8, -15, -7, -9, 2, -7, -19, -3, -8, -4, 5, -12, 10, -15, 18, 1, -23, 23, -15, -6, 2, -9, 6, -32, -21, -9, 1, -34, -25, -15, 0, -14, -13, -13, 30, 4, -4, 0, 13, 5, -3, -18, -41, 21, 19, 1, -13, -6, 4, 3, -4, -11, -4, -7, -17, -2, -4, 3, 2, 9, 6, -4, -8, 2, -4, 15, -15, -6, 6, -5, -8, -14, -13, -18, -5, -4, -6, -18, 7, -9, 1, -1, 4, 9, -22, -7, 7, 3, 1, -12, -15, 16, 8, -7, -13, -7, -2, 7, 18, -9, 11, 8, 3, 1, -4, 16, 7, 2, -6, 7, 7, 1, -7, 1, -3, 7, -1, 8, 0, 4, -3, -10, -10, -11, 4, -5, 5, -1, -3, -9, 4, -9, -8, -9, 3, -7, -1, 8, -4, 7, 0),
    (12, -7, 4, -7, -15, 7, -6, -15, 13, -9, 11, 16, -26, 1, 5, -5, -7, 17, -11, -6, 5, -17, -3, 1, 3, 11, 3, 10, 20, 8, -1, 13, -8, -10, -9, -5, 23, 6, 12, -1, -10, 2, -30, -11, 2, 2, -12, -18, 46, -23, 16, -7, -19, 5, -16, -42, 11, -21, 16, 17, -22, 7, 10, 15, -15, -27, -7, 22, 9, -21, -15, 13, 7, 14, 11, 25, 48, 14, -4, 31, -39, 59, -12, 2, 21, 1, -13, -3, -16, -35, -51, -25, -11, -5, -24, 3, 26, -9, 18, 3, -21, 2, -13, -36, 10, -23, 2, 1, -4, 2, 3, 16, -25, -20, 0, 32, 20, -27, -19, 3, 22, -10, 5, 46, 41, 4, 0, 20, -23, 54, -7, 3, 23, 13, -22, -1, -16, -37, -25, -21, -21, -17, -20, 0, 13, -6, 14, 7, -4, 10, 5, -22, 4, 9, 6, 3, 11, 5, 3, 9, 0, -14, -14, 16, 18, -15, -14, 5, 9, -11, -2, 45, 18, -7, 4, -4, -10, 40, 5, 5, 3, 7, -13, 3, -1, -26, 5, -9, -17, -21, -7, 8, 16, -27, 18, -15, -19, 13, -26, -40, 13, 7, -20, 14, 3, 8, -15, 7, 9, 2, -34, -17, 12, -6, -23, -20, 4, 17, 3, -6, 11, 6, 2, 4, -17, 5, -4, 4, 22, -14, 7, 16, 2, -23, -16, -23, -5, 2, -5, -9, 27, -19, 9, -1, -34, 7, -51, -57, 19, 6, -5, 3, 14, 10, -19, 32, -19, -47, -24, -33, 15, -21, -35, -19, 3, 26, 0, -22, 35, 22, 13, 14, -35, 28, 1, -5, 35, -8, -10, 21, -9, -46, -11, -36, -26, -4, -9, -29, 23, -13, 15, -2, 2, 0, -40, -35, 15, 6, -6, -12, 8, -7, -24, 22, -30, -23, -29, -17, 21, -22, -23, 8, 20, 7, -12, -1, 30, 26, 14, 15, -26, 25, 1, -1, 45, 4, -16, 12, 13, -42, -19, -35, -30, -12, -19, 2, 9, 0, 22, -8, 13, -9, 9, -18, 13, -14, 2, -7, 1, -18, -4, 5, -2, -12, -8, 12, 17, -17, -12, 4, 9, -5, 7, 1, 15, 4, 7, 9, -6, 13, 15, 18, 16, -4, -18, 22, 2, -14, -20, -19, -14, -21, -3, 5, 2, 2, 29, -8, -5, 3, -12, -12, 1, -1, 2, -3, 5, 14, -4, 1, 6, -16, -14, 4, 6, 1, -5, -12, -2, 5, 11, -9, 8, 6, -1, -2, -26, -11, 16, -4, 9, -22, -13, 7, 5, -7, -3, -2, -9, 10, 11, -10, 10, -20, 30, 5, -15, 0, -6, -15, -2, 7, 2, 15, 8, 11, -5, 16, -15, -23, -39, -11, -9, -10, -19, -29, 8, 19, 11, -22, -4, 13, -12, 10, -27, -10, 11, 5, 18, -23, -17, 5, 6, -8, 7, -14, -14, 2, -9, -17, 14, -8, 19, 1, 2, -5, -5, -1, 4, 17, 9, 15, 8, 1, -19, 5, 5, -14, -40, 2, -4, -11, 11, -17, 2, -7, -6, -9, 4, -7, -13, 11, -18, -2, 8, 0, 15, -7, -9, 9, 19, 2, -10, -11, -1, -10, 1, 2, 9, -14, 0, -1, -3, -13, 1, 4, 2, 5, 15, 1, 18, 4, -3, -2, -12, -3, -16, 6, 5, -4, 1, -8, -4, -16, 1, -2, 4, 0, -18, 0, -1, -4, 8, -1, 5, 0, 11, 18, -3, 11, 2, -2, 5, 1, 12, 5, 8, -8, 28, -8, -12, 4, -4, -2, 6, 12, -3, -7, 2, 6, 9, -6, -7, 5, -15, 10, 0, -11, -5, -9, 6, 1, 9, -9, 1, 2, -8, 2, 8, 6, 18, -1, -4, -16, -9, 11, 6, -4, 6, 8, -13, 2, -1, 5, -5, -19, 14, -1, 1, 9, -3, 2, -10, 17, -1, -1, 3, -5, 6, -8, 1, 0, -20, -11, -6, 14, 2, 8, 6, -5, 23, 1, -5, -3, -15, -3, -6, -4, 11, 4, 4, -16, -20, -6, 3, 3, 7, 14, -6, 10, -1, 0, -8, -15, -1, -2, 4, 5, -8, 5, -15, -4, -4, 6, 11, -7, -1, -3, -13, -2, 0, 2, -4, -1, 10, 4, -9, -4, 9, -4, 9, 5, -6, -17, 3, 5, -12, -7, 3, -11, 7, -28, 9, -5, 9, 17, 11, 11, 13, -8, 11, -7, -12, -24, 5, -15, -7, -8, -5, 3, 4, 5, 4, -3, 7, -11, -13, 7, -6, -14, 2, 0, -12, -5, -7, 9, -11, -9, 16, 8, -9, 5, -17, 14, 4, 5, -14, -10, -15, 9, -12, -4, -10, -3, 8, 10, -2, 2, 1),
    (-33, 19, -25, 19, -30, -22, -16, 6, -2, -13, 7, 26, -13, -6, -20, 13, 21, 6, -30, -10, -9, -52, -34, -2, -25, 30, -38, 22, 30, -2, -9, -10, 23, -3, -20, -29, 4, 14, -7, 17, -17, -15, -10, -18, -8, 9, -21, -15, -40, -4, 9, 16, -6, -29, -30, -5, 20, -13, 2, 14, -42, 11, 6, 23, 8, -18, -55, 3, -12, -50, -41, 21, -1, 35, -36, 31, 25, -8, -23, -23, 10, 29, -27, -38, 4, 17, -13, 4, -33, -60, -44, -33, -1, -6, -30, -4, -49, -1, -1, 8, -19, -23, -25, -17, 12, -11, -4, 15, -35, 1, -10, -11, -25, -13, -21, 7, 5, -34, -23, 4, 14, 1, -21, 36, 14, 11, -13, -2, -13, 16, -19, -27, -10, -11, -24, 14, 4, -26, -30, -30, -4, -1, -28, -7, -9, -12, 3, 4, -38, -13, -19, -19, 10, -15, -12, 17, 1, -9, 10, 3, -16, 3, -11, -8, 2, -25, -5, 9, -11, -15, -12, 20, 15, 10, -12, 9, 5, 5, -13, 6, 6, 4, -8, 0, 0, -9, -25, -19, -5, -4, -13, -3, -18, 26, -24, 26, -6, -14, -34, 18, -6, -4, 30, 26, 2, 18, 24, 23, 19, -2, -10, 9, -21, -42, -18, 21, -20, 18, -29, 31, 11, 25, -18, 1, 18, -3, -33, -12, -4, 13, 8, 9, -14, -20, -10, 23, 17, -6, -4, 12, -9, -3, -10, 14, -6, -6, -53, -10, 9, 14, 17, 15, -9, 0, 24, 18, 19, -9, -31, 25, -22, -51, -32, 20, -21, 22, -35, 17, 31, 14, -30, 4, 9, 8, -27, 1, 13, 31, -1, 24, -36, -45, -10, 30, 15, -11, -8, 5, -6, -12, -11, 6, -34, 7, -30, -21, -3, 13, 19, 18, -10, 1, -8, 11, -29, -10, -39, 20, 2, -32, -21, 15, 1, 15, -31, 20, 14, 31, -26, 11, -1, 11, -7, -2, 14, 7, -15, 13, -33, -27, -20, 24, 13, -10, -13, 2, -2, -3, -10, -7, -17, 2, -10, -7, 2, 0, -4, -2, -7, 1, -15, -17, -9, -5, -8, -5, 9, -10, -20, 0, 1, -3, -11, 10, 10, 0, 0, 8, 8, 6, -3, -10, 4, -1, -11, -1, -4, -1, -24, 7, -11, -4, 19, -18, -8, -1, -11, -11, -6, -6, 16, 19, 0, 4, 24, 9, 16, 21, 15, 3, -6, 18, -14, 7, 12, -53, 0, 24, -19, 24, -28, 24, -8, 18, -9, -1, 32, -13, -21, 23, -9, 6, 13, -3, -20, 8, -25, 20, 14, -18, 5, 1, 6, -22, -6, -6, -8, 1, -1, 9, 4, 7, 29, 3, 0, 9, 14, -10, 15, 24, -24, 16, 16, -46, -18, 5, -14, 38, -23, 7, 0, 23, -38, 0, 14, -16, -12, 24, -8, 9, 7, 2, -49, 5, -14, 21, 40, -19, 4, 15, -1, -16, 1, -7, -8, 6, 1, 0, 2, 8, 24, 19, -5, -10, 12, -13, -25, 17, -43, 31, -3, -28, -11, -6, -20, -8, -13, 17, -15, 13, -38, 15, 18, 1, -1, 11, -1, 6, -1, -6, -68, -17, -30, 27, 20, -6, -3, 15, 2, -15, -4, -15, -26, 4, 8, 8, 8, 5, 2, 4, 12, -14, 9, -5, -6, 19, -17, 11, -18, 6, -14, 7, -25, 0, 3, -3, -15, 0, -29, -3, 7, 11, -1, -1, -4, 7, 18, -5, -17, 3, -12, 20, -7, 30, 8, -1, 6, -32, -4, -8, -15, 0, 5, -2, 24, 7, 10, 9, -13, 16, 13, -4, -22, -2, -20, 0, -2, 15, -7, 3, -36, -14, 4, 11, -10, 21, -26, 11, -5, -25, -13, 11, -6, 1, 12, -7, -38, 0, -33, 11, 0, 0, 3, -6, -4, -27, 13, -21, -8, 12, 5, 9, 14, 2, 21, 3, -20, 1, 11, -15, 0, 22, -31, 9, -6, -14, -2, -7, -31, -9, -3, 2, -8, 18, -32, 1, -8, -15, -3, 9, -3, 12, 13, -7, -25, -6, -19, 18, 6, 4, -2, -2, -1, -18, 12, -7, -9, 10, -7, -2, 22, 12, 19, -9, -12, -9, -1, -11, -16, -3, -7, 10, 8, -14, 7, -5, -28, 0, 9, 0, -17, 3, -26, 5, -4, -7, 9, 8, -10, -2, 7, 10, -20, -17, -15, -8, -4, 11, -1, 1, -6, -20, 7, -1, -13, 2, 11, -9, 12, -5, 6, 12, -25, -1, 5, -18, -6, -15, -10, 7, -3, -13, 3, 3, -7, 6, -14, 23, 12, -7, -2, -6, -11, -4, 2, -6, 1, -2, -7, 20, -21, 3, -7, 3, -3, -22, 11, 4, -13),
    (-17, -4, 2, -13, -2, -11, 13, 18, -41, 25, 3, -5, 28, 5, 2, -12, -22, -32, 42, -3, -18, 26, 10, -19, 17, -37, 10, -4, -11, -27, -6, -47, -24, -1, 10, 11, 0, -5, -21, -1, 21, 2, 27, -10, -18, -34, 2, 9, -53, 15, -8, -20, 24, -24, 8, 18, -23, 8, 1, 11, 21, 8, -1, -10, -31, -4, 36, -20, -13, 5, 21, -17, 19, -51, 7, -1, -8, -34, 11, -39, -14, -11, 19, 18, -14, 2, 5, 1, 37, 20, 31, 2, -17, -18, 21, 21, -50, 1, -9, -12, -1, -15, 8, 12, -26, 7, -1, -9, 18, -7, 0, -3, -7, 1, 24, 1, 0, -6, 19, -23, 13, -10, 14, -26, -21, -24, 12, -38, -10, -20, 16, 9, -2, 6, 14, -7, 32, 7, 30, 18, -9, -8, 14, 27, -12, 2, -1, -6, -17, -13, 7, 2, -22, -10, -6, -8, 8, -5, 4, -9, 0, 8, 1, -13, -13, 6, 6, -4, -1, -9, 1, -29, -10, 0, 3, -24, 1, -15, 11, 9, -3, -11, -8, 2, -7, 19, -5, 12, -9, -1, 0, 3, -6, 30, 6, -5, -18, -21, 12, 11, -26, 15, -21, -33, 7, -23, -19, -9, -20, -8, 29, -32, -9, 18, 15, -11, 7, -42, -1, -30, -22, -27, 27, -44, -16, -1, 12, 9, -28, 17, -13, 7, 22, 21, 12, -18, -32, -21, 4, 3, -33, 40, -16, -18, -11, -26, 25, 28, -8, 3, -2, -16, 15, -11, -14, -14, -29, 5, 43, -39, -13, 16, 30, -10, 4, -45, 1, -9, -6, -44, 41, -34, 9, -9, 3, 28, -18, 29, 5, -4, 31, 36, 19, -19, -24, -5, 16, -7, -38, 20, -15, -10, -9, -28, 27, 16, -10, -2, 15, -15, 12, -9, -9, -16, -9, 0, 31, -34, -19, 9, 16, -21, -7, -8, 9, -24, 0, -23, 32, -34, 11, -3, 3, 14, 5, 10, 11, -17, 34, 32, 20, -6, -7, -4, 11, 4, -25, 1, -16, -4, -14, -13, -6, 9, -3, -8, 9, 10, 2, 0, 3, -5, 2, 2, 7, -6, -5, -2, 9, -4, 0, -6, 11, -14, -6, -13, 1, -8, -4, -10, 9, -3, -5, -4, 10, -3, 8, 23, 5, 10, -3, 12, 12, 15, -14, 12, -25, 13, -12, -4, -28, -24, -27, -1, -8, -2, 5, -25, -35, 4, -10, -28, 25, -32, -14, 12, 9, -10, 14, -31, 2, -35, -7, -14, 25, -25, -29, 8, 9, -37, -18, 14, -16, -18, 17, 13, 9, -16, -30, -5, -17, -4, -21, 25, -31, 12, -25, -19, 7, -15, 14, -1, -19, -14, 1, -10, -25, 7, -35, -36, 30, -18, -13, 29, 11, -22, -1, -53, 6, -16, -6, -42, 33, -22, 1, 1, -9, 1, -7, 11, -5, -29, 37, 11, 13, -20, -45, -11, -27, -7, -7, 17, -27, 8, -10, -25, 5, -1, 13, -3, 2, -24, 5, 9, -4, -12, -32, -22, 29, -14, 0, 10, 9, 0, 15, -2, -8, -13, 4, -13, 25, -15, 2, 2, -9, -7, 12, 11, -4, -25, 22, 20, 13, -18, -9, 5, -18, 2, -15, -1, -20, -10, -3, -11, 10, 8, -11, -6, -7, 1, -13, 10, 0, -16, -17, -5, -5, -8, -6, 11, -1, -17, 3, -3, -13, -5, -9, -3, 6, -11, -12, -3, -15, -7, 5, 9, 7, -9, 0, 14, 2, 0, -9, -25, -13, 12, 2, 18, -31, 7, -6, -1, 5, -11, -38, -35, -11, -7, 1, 0, -9, -2, 1, -3, 18, -7, -6, 1, 7, 0, 5, 4, -9, -7, -5, -5, 3, -41, -7, 13, -9, -14, -5, -9, -23, -28, 13, 8, 11, -12, 0, -4, -12, 3, -3, 19, -45, 47, -8, 2, 12, -10, -42, -22, -8, -24, 3, 16, -22, 14, -39, -22, 20, -13, 9, 9, -9, 1, 32, -2, -11, -6, 3, -15, 22, -26, 14, 11, -7, -44, 4, 10, -28, -16, 17, 9, 16, -7, -4, -26, -15, -9, -9, 11, -34, 12, 4, -6, 3, -10, -32, -27, -7, -26, 10, 13, 4, -13, -11, -3, 7, -6, -13, 0, 5, -10, 19, 6, -2, -12, -2, -3, 15, -9, -9, -1, -1, -15, 8, 4, 1, -17, 10, 17, 14, -17, -2, -8, -13, -7, -1, -5, -27, 7, 4, 0, 8, -2, -28, -14, 4, -8, 15, 0, 1, -2, -23, -1, 8, -13, -3, 3, 0, 6, 6, 4, -3, -31, 10, 2, -13, -14, -6, -13, 3, -3, -6, -6, -1, -19, 20, 4, 2, 2, 9, -6, 3, 6, -1),
    (3, -9, -11, -6, -2, 1, 7, -26, 3, -17, -7, -9, -6, 2, -9, -20, -8, 10, -1, -29, 21, 6, 1, 8, -11, 15, 4, -23, 8, 28, 9, 20, -2, 0, -13, 18, -6, 17, 17, -34, -6, 11, -26, 3, -2, 23, -10, 10, 18, -12, -13, 3, -9, 4, 16, -20, -1, -13, -1, -17, 1, 1, -16, -24, 1, 7, 4, -35, 10, -1, 5, 2, -31, 6, 8, -24, 4, 22, 7, 28, 1, 2, -1, 28, -9, 14, 4, -15, -16, 11, -16, 15, -2, 26, -4, 14, 24, -11, -6, 7, 7, -1, 11, -11, -4, -10, 3, -12, 0, 7, -14, -10, -2, -1, 8, -25, -8, -11, 11, 1, -13, 3, 11, -4, -3, 13, 0, 15, 10, 10, -14, 13, -10, 15, 6, -5, -16, 9, -3, 11, -2, 17, 0, 6, 8, -13, 8, 10, 10, 0, -8, -6, 15, 7, -4, -10, 0, -5, -14, -4, 3, -7, 2, -16, 15, -8, 9, -5, -12, 10, 7, 3, -6, 12, 8, 10, 12, -1, 7, 11, -2, 9, 9, 3, -9, 0, -3, 6, -1, -4, 0, 5, -2, -22, -29, 10, 17, 15, -2, -44, -2, -39, 12, -15, -14, 0, -19, -1, 2, 8, -5, -14, 17, 15, -9, -3, -4, 20, 2, -22, -22, 15, -1, 11, 1, 21, -5, 27, -22, 4, 13, -33, -11, -1, -14, 2, 0, 14, -32, -15, 10, -29, -13, 7, 14, 17, 16, -33, -6, -20, 13, -28, -14, 5, -19, -21, -5, 5, -3, -29, 18, 3, -14, 3, -28, 28, 2, -23, -17, 3, 13, 14, -1, 17, -13, 21, -20, 13, 3, -34, -14, 16, -18, -6, -14, 15, -34, -50, 26, -22, -2, -1, 7, 8, 15, -19, -3, -17, -4, -18, -3, 15, -12, -12, 3, 12, 1, -24, 1, 0, -19, 16, -17, 21, -3, -11, -13, 18, 6, 11, 2, 16, -11, 23, -10, -8, 0, -19, -13, 8, -32, -4, -5, 24, -28, -36, 12, -5, -4, -3, 8, -1, 2, -16, 5, 3, 10, 6, 7, -1, -4, -2, 8, -10, 2, 10, -2, 0, -5, 8, -12, 14, 1, 5, 2, 2, -2, 13, 10, 11, 1, 13, -8, 1, 5, -15, 13, 0, -13, 5, 10, 8, -17, -14, 3, -17, -18, 29, 3, 16, 13, -21, -12, -5, 20, -13, -10, -3, -10, -12, -12, -2, 5, -7, 4, 28, -8, 1, -13, 6, -6, -21, -11, 8, -7, 15, 2, 28, -4, 0, -12, 13, 10, -12, -19, 0, -3, 10, 1, 11, 18, -15, 15, -33, -2, 21, 22, 16, 14, -19, -19, -14, 16, -41, -6, -3, -11, -13, -11, -9, -5, -13, 6, 17, -22, -5, -15, 26, -19, -19, -19, 10, -7, 11, 14, 12, -2, -1, -24, 13, 15, -14, -23, -2, -10, -2, -4, 4, -4, -27, 24, -23, -2, 8, 26, 5, 7, -13, -1, 0, -1, -21, -13, 3, 1, -3, 11, -15, 0, -11, 2, 5, -23, -1, -11, 16, -16, -10, -17, 27, -12, 18, 3, 3, -4, 1, -16, 0, 0, 0, -29, 9, -33, 4, -3, 15, -1, -12, 10, 6, -7, -3, 18, 0, 6, -8, -11, -9, 7, -9, -22, -4, 1, 14, 1, -8, 2, -4, 6, 1, -10, -7, 6, 1, -21, -8, -13, 10, 0, 19, -1, 10, 1, -8, 0, 1, -18, 18, -12, 9, -13, 8, 3, -1, 6, -1, 2, -1, 6, 9, 16, 6, 1, 14, 3, 7, 5, 0, 0, 9, -6, 1, -1, -5, -1, 1, 6, 1, 9, -2, -18, 2, -11, 10, 1, 14, 11, 11, 10, 9, 1, 10, -15, 16, 3, 16, -22, 16, 4, -1, -3, 5, 9, -3, 19, -12, 3, 11, 12, 13, 6, 7, 1, 12, 14, 6, 7, -9, 7, 1, 19, -11, -9, 2, 11, 6, -13, 8, -15, 10, -16, 8, 5, 14, -10, 11, 7, -8, 13, 9, 7, 13, -9, 17, -7, -1, 5, 14, -6, 1, 17, -15, 8, 5, -4, 8, 9, 6, 2, 9, -6, 12, 7, 5, -4, 1, -7, 3, 24, -3, 1, 9, -5, -6, -4, -10, -13, 6, -1, -15, -17, 7, -4, -6, -8, -11, -1, 7, -7, 13, -7, 0, 2, 14, -15, -12, 0, 2, -10, 0, 11, 12, -11, -18, 2, -2, 2, 5, 1, -6, -12, -14, -3, -18, -1, -16, -3, -6, 14, -15, -7, 8, 4, 0, -5, -6, 2, -16, 3, -2, 3, -2, -1, 7, 15, 7, 3, 6, -2, -12, -10, 0, -4, -5, 3, 28, -12, -7, 7),
    (33, -2, -20, 12, 10, -4, -11, -22, 9, 8, 1, -8, 10, 3, 14, -14, -8, 1, 22, 23, 11, 24, 10, -2, -21, -14, -22, -11, 18, 31, 6, 5, -1, 9, -16, 1, -12, 14, -5, -11, -25, 15, -12, 12, 7, 1, 16, 19, 51, -12, -13, 3, -8, -11, -4, -20, 4, 10, 16, -14, 11, -1, -7, -4, -28, 3, 11, 34, 9, 12, 4, -11, -21, -18, -7, -36, 16, 39, 21, 18, -5, -7, -11, 2, -7, 18, -10, 3, -32, 22, 6, 31, 17, 4, 16, 24, 30, -4, -1, 9, 1, -11, -9, -22, 16, 32, 5, -24, 16, 0, -17, -15, -15, -2, -8, 3, -4, -3, 9, -6, -14, -15, 2, -44, 0, 31, 11, 9, -13, -14, -8, 12, -4, 18, -2, 4, -39, 16, 6, 25, 10, 13, 10, 21, 13, 10, 12, -8, -8, 11, 6, -11, 1, 17, -1, -27, 1, 1, -3, -16, -8, 1, -2, -2, 5, 10, 6, -21, -9, -2, 21, -17, -11, 4, -1, 2, -13, -14, 0, 3, -2, 13, -5, 21, -19, 9, -10, 19, -8, 3, 10, 5, 26, 11, -20, -31, -2, -7, -34, -9, 26, 6, -49, 13, -5, -11, 3, 4, -22, -4, 28, 21, 11, 18, 14, -13, -11, -3, 1, 11, 12, 28, 5, 2, -21, 11, -2, -8, 1, -9, -3, 8, -14, 0, 12, 3, 26, 2, -11, 18, 18, 28, -13, -22, 6, -7, -34, -15, 27, 3, -56, -25, 11, -11, -11, 18, -50, 7, 20, 16, -1, 17, 9, -32, -15, -17, 5, -21, 17, 30, 27, 13, -25, -17, -12, -9, 5, -6, -12, 8, -23, 14, 18, 9, 48, -5, -25, 30, 6, 21, -5, -15, 13, -14, -32, -12, 13, 11, -42, -28, 18, 9, -5, -1, -17, 8, -4, 0, -15, 20, 4, -15, -18, -20, 5, -36, 15, 18, 16, 9, -24, -14, -8, 5, 15, 11, -5, 4, -20, 13, 27, 5, 27, 1, -16, 24, -1, 13, 10, -1, 0, -2, -13, 1, -7, -4, -6, 8, 10, -10, 9, 0, -3, 7, -9, 5, -3, 13, -4, -7, -5, 8, 17, -20, -12, 8, -5, 0, -17, -13, 7, 8, -6, 8, 9, 10, -6, 13, -5, 18, 4, 7, 1, 7, 4, 21, -7, -28, 6, -10, -33, -23, 24, 10, -22, -4, 9, -16, -3, 5, -11, -10, 11, -9, -12, 30, 23, -9, -1, -3, 6, 9, 6, 0, 10, 10, -45, -10, 9, -13, 13, 4, 6, 5, 6, 5, 7, 0, -16, 10, -16, 1, 6, 32, -15, -5, 4, -12, -33, -18, 40, 7, -43, -31, 4, -19, -15, 11, -38, -13, 10, -10, -30, 21, 26, -22, 7, -41, 7, -22, -9, -1, 18, 3, -44, -21, 4, -6, 10, -6, 7, -10, 8, -12, 26, 22, -16, 12, -34, 0, 5, 18, -11, -1, -11, -15, -27, -17, 18, 2, -38, -28, -1, 1, -2, -4, -26, -10, 9, -4, -24, 24, 2, -14, 23, -7, 6, -15, -16, -11, 20, -5, -42, -23, -14, -7, 3, 3, 12, -28, 13, 1, 12, -1, -7, 18, -30, 6, -10, -5, -2, -14, 1, -1, 4, -9, 0, -1, -8, 1, -24, -10, 7, -2, -10, 1, -3, 1, 3, 12, -6, 9, 5, -3, -19, -6, -2, 11, 3, -17, -14, -33, -6, 0, 1, 11, 4, -12, -2, 7, 1, -12, -16, -12, -12, -6, -4, -3, -18, 7, -15, 2, -14, -14, -36, -2, -15, -9, 2, 4, -14, 1, -11, 2, 0, -15, 3, 8, 3, 6, 12, 17, 6, -1, 3, 1, 5, -15, -18, -1, -5, -4, -6, -10, -9, -8, 8, 2, 17, -2, -6, -22, -6, -2, -9, 6, -38, 25, -18, 7, -14, -15, -16, 2, -11, -20, 8, -6, -14, 0, -23, -19, 23, -22, 4, 14, 6, -4, 21, 3, 12, -13, -12, -12, 11, -27, 0, -9, 6, -17, -1, -17, -4, -19, 14, -1, 16, -19, -14, -32, -20, -6, -4, -2, -29, 3, -9, -4, -18, -15, -30, -11, -15, -13, 4, 15, -13, 2, -5, -11, -4, -3, -5, 0, -7, -5, 12, 6, 2, 2, -8, 10, -1, -3, 9, -9, 10, -19, 1, -1, -2, -17, 1, 7, 19, -2, 5, -24, -20, -4, 13, -3, 4, 7, -6, -16, 1, -7, 8, 10, -13, 7, 18, -14, 2, 0, -15, -5, 4, 1, 0, 10, -3, -6, -10, 10, 9, -6, -1, -3, -9, 15, -18, -12, 12, -5, -2, -1, -5, -2, -12, -8, -12, -11, -11, 5, -3, -9, -6)
  );
  ----------------
END PACKAGE CNN_Data_Package;
