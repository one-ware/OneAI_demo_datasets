library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.numeric_std.all;
use work.CNN_Config_Package.all;

PACKAGE CNN_Data_Package is
  CONSTANT Layer_1_Columns    : NATURAL := 128;
  CONSTANT Layer_1_Rows       : NATURAL := 128;
  CONSTANT Layer_1_Strides    : NATURAL := 1;
  CONSTANT Layer_1_Activation : Activation_T := relu;
  CONSTANT Layer_1_Padding    : Padding_T := same;
  CONSTANT Layer_1_Values     : NATURAL := 1;
  CONSTANT Layer_1_Filter_X   : NATURAL := 3;
  CONSTANT Layer_1_Filter_Y   : NATURAL := 3;
  CONSTANT Layer_1_Filters    : NATURAL := 8;
  CONSTANT Layer_1_Inputs     : NATURAL := 10;
  CONSTANT Layer_1_Out_Offset : INTEGER := 3;
  CONSTANT Layer_1_Offset     : INTEGER := 1;
  CONSTANT Layer_1 : CNN_Weights_T(0 to Layer_1_Filters-1, 0 to Layer_1_Inputs-1) :=
  (
    (52, 19, 20, 10, -30, 15, 26, -5, 51, 2),
    (-31, -25, -51, -17, -25, -17, -50, -27, -32, -2),
    (-9, 23, 39, 3, -42, 56, -48, -37, 6, 0),
    (-13, 0, 26, 28, 9, 10, 50, -9, 69, 2),
    (19, 31, 35, -23, -4, -6, -32, -66, -38, -1),
    (27, 34, 7, 30, -6, -25, -12, -29, -57, -1),
    (26, 46, 10, 37, 36, -7, 14, -3, -14, -1),
    (71, -60, 36, -43, -39, -15, -62, 19, 16, -1)
  );
  ----------------
  CONSTANT Pooling_1_Columns      : NATURAL := 128;
  CONSTANT Pooling_1_Rows         : NATURAL := 128;
  CONSTANT Pooling_1_Values       : NATURAL := 8;
  CONSTANT Pooling_1_Filter_X     : NATURAL := 2;
  CONSTANT Pooling_1_Filter_Y     : NATURAL := 2;
  CONSTANT Pooling_1_Strides      : NATURAL := 2;
  CONSTANT Pooling_1_Padding      : Padding_T := valid;
  ----------------
  CONSTANT Layer_2_Columns    : NATURAL := 64;
  CONSTANT Layer_2_Rows       : NATURAL := 64;
  CONSTANT Layer_2_Strides    : NATURAL := 2;
  CONSTANT Layer_2_Activation : Activation_T := relu;
  CONSTANT Layer_2_Padding    : Padding_T := same;
  CONSTANT Layer_2_Values     : NATURAL := 8;
  CONSTANT Layer_2_Filter_X   : NATURAL := 3;
  CONSTANT Layer_2_Filter_Y   : NATURAL := 3;
  CONSTANT Layer_2_Filters    : NATURAL := 12;
  CONSTANT Layer_2_Inputs     : NATURAL := 73;
  CONSTANT Layer_2_Out_Offset : INTEGER := 4;
  CONSTANT Layer_2_Offset     : INTEGER := 0;
  CONSTANT Layer_2 : CNN_Weights_T(0 to Layer_2_Filters-1, 0 to Layer_2_Inputs-1) :=
  (
    (-39, -10, 22, -11, 32, -5, -9, 34, -6, -50, 60, -3, 29, -9, -6, 29, 40, -16, 10, 11, -12, -68, -12, -18, -11, 14, -49, 4, 20, 15, -4, 28, -21, -38, 9, 19, -24, 29, -20, 68, -8, -34, 8, 3, 12, 13, 3, 52, -3, 9, -37, 29, -46, 13, 9, 30, 23, -31, -9, -23, -40, 37, -9, 36, -46, 23, 2, -28, 29, 35, 28, 59, -3),
    (-23, 8, -17, -16, 8, 37, 13, 41, -11, -2, -1, 31, -1, 50, 44, 42, 41, -62, -3, 43, 7, -10, 15, 4, -35, 16, -19, -4, 43, 48, 24, 30, -37, 20, -13, -8, 63, 69, 42, 32, -18, -39, -12, 2, 26, 31, 42, -8, -20, 13, -36, 8, 39, 30, -9, -28, -31, 29, -29, -19, 51, 64, -15, -11, -5, -20, -22, -5, 1, 40, -28, -9, -4),
    (16, -33, -22, 45, -74, -58, 5, -37, 20, -8, -12, 18, -1, -93, -3, -42, 30, 9, -19, 7, -30, -34, -13, 10, 45, -69, 1, 1, 12, -21, 19, -13, -30, -66, 13, 36, 22, -65, -7, -43, 35, -54, 4, 23, 7, -59, -34, -23, 35, -13, 14, -10, -4, -18, 26, 12, -15, -35, 7, 24, 17, -24, -30, -5, -9, 55, 8, 3, 32, -12, 4, 12, -1),
    (-25, 49, 27, -42, -21, 5, 28, 0, -5, 52, -61, -42, 5, -48, -31, 6, -8, 5, -25, -3, -33, 3, -45, 10, -11, 30, -45, -5, 6, -81, -18, -30, 13, 16, -27, -3, 40, -30, -8, -34, -12, -6, -35, -32, -15, -25, -17, 4, 18, -34, 7, 42, 98, 4, -9, 15, -3, 5, 28, 10, 53, 2, -12, 29, 12, -12, 10, 7, 16, -7, -20, 25, -3),
    (-16, 14, 29, -19, 3, 5, 16, 5, 11, -51, 16, -3, -33, 1, 40, 14, 28, -43, 17, -6, 3, -3, 38, 7, -5, -4, 19, -15, 14, 10, -4, 24, -18, -91, 32, 4, 5, 16, 21, 47, 24, -9, 22, 10, 0, -18, 30, 25, -63, 58, -16, -37, 12, 46, -46, 5, -16, -20, 27, 12, 20, 30, -8, 6, 3, -14, 44, 14, -32, 1, 17, 11, -10),
    (-37, 25, -35, 1, -35, -87, -24, -33, -44, 42, -42, 15, -34, -72, -14, -30, -65, -27, -30, -38, -15, -72, -68, 13, -11, -10, 24, 20, 23, -4, 37, 29, 14, -49, 51, 15, 41, -49, 42, 13, 2, -8, 32, 1, 52, -43, 10, 28, 16, 24, 21, -23, 15, 16, 5, 31, -14, 13, 43, -11, 12, -14, 36, 21, -20, -8, 28, 3, 12, -6, 1, 4, -4),
    (-29, -10, 27, -12, 27, -17, 5, 30, -23, -6, 47, -2, 58, 16, -7, 35, 2, -2, 62, 0, 47, 30, 17, 35, -4, 16, -45, 11, 22, -35, 1, -54, -4, 62, -20, -16, 42, -9, -39, -23, 10, -24, -12, -26, 27, -23, -18, -19, 31, -11, -6, 21, -37, -36, 26, -41, -4, 49, -26, 26, -10, -40, 12, -47, 5, 26, -32, 14, -25, 9, -12, -47, -2),
    (16, 14, -10, -9, 45, 7, -23, -25, -27, 29, -25, -4, 58, -47, -22, -45, -36, 17, 34, -4, 30, -38, -12, -14, -10, 11, 18, 54, -29, -25, 25, -29, -5, -11, 3, -7, -82, -36, -11, -47, -24, 48, 1, -53, -14, -35, 2, -19, 1, -14, 14, 41, -52, -27, 43, -12, 44, -14, 40, 33, -55, -26, 14, -34, -3, 8, 29, -27, -65, -59, 0, 5, -3),
    (-28, 38, -24, -13, -40, -14, -74, -5, 2, 49, 1, 11, -70, -5, -39, 3, 9, -21, 44, 5, -38, 40, -17, 36, -43, 45, -10, -33, -42, -17, -61, -14, -33, 32, 14, 22, -68, 10, -5, 14, 10, -10, 28, 38, -19, 44, 36, 85, 0, 11, 15, -21, -10, -26, -44, -9, -4, -23, 30, 28, -34, -5, 19, 34, 36, -2, 4, 44, -28, 16, 37, 64, 3),
    (22, -42, 7, 20, 8, -14, 14, -2, -23, -50, 8, 10, -25, 2, 28, -17, 25, 7, -2, 0, -7, -27, 2, -44, -4, -63, -1, 24, 2, -9, 36, -15, 1, -122, 7, 7, -36, -35, 9, -41, 18, 5, 30, -4, -21, -44, 8, -37, 10, -37, -19, 20, -29, 2, 13, -4, -23, -5, -6, 36, -31, -27, 26, 7, 41, 8, -5, 34, -17, -77, 5, -9, -9),
    (21, -16, -9, 15, -28, 28, 43, 35, -1, -98, 0, 13, -51, 20, 33, 34, 8, -30, 19, -12, -25, 20, 26, 4, 20, -65, 7, 6, -45, 10, 43, 29, -54, -103, 47, 8, -42, 29, 44, 17, -23, -58, 30, 4, -20, 14, 8, -8, 19, -62, 17, -11, -26, -8, 25, 5, -3, -60, 28, -10, -19, -18, 25, 15, -11, -39, 23, 33, 6, 4, 2, 15, -4),
    (20, -49, 26, -25, 12, -28, -22, -6, 31, -105, 36, -11, 32, -52, 27, -12, 4, 6, 4, 28, -7, -46, 27, -25, -38, 31, 34, -31, 62, -9, 4, 21, -2, 2, 42, -4, 66, -9, -14, -15, 14, -10, 41, 1, 77, -8, 9, 4, 26, 1, -61, 23, 37, -71, -28, -39, -19, 8, -29, -12, 62, -40, -43, -35, 0, -1, -4, -9, 71, -35, -6, -8, -5)
  );
  ----------------
  CONSTANT Layer_3_Columns    : NATURAL := 32;
  CONSTANT Layer_3_Rows       : NATURAL := 32;
  CONSTANT Layer_3_Strides    : NATURAL := 2;
  CONSTANT Layer_3_Activation : Activation_T := relu;
  CONSTANT Layer_3_Padding    : Padding_T := same;
  CONSTANT Layer_3_Values     : NATURAL := 12;
  CONSTANT Layer_3_Filter_X   : NATURAL := 3;
  CONSTANT Layer_3_Filter_Y   : NATURAL := 3;
  CONSTANT Layer_3_Filters    : NATURAL := 16;
  CONSTANT Layer_3_Inputs     : NATURAL := 109;
  CONSTANT Layer_3_Out_Offset : INTEGER := 5;
  CONSTANT Layer_3_Offset     : INTEGER := 0;
  CONSTANT Layer_3 : CNN_Weights_T(0 to Layer_3_Filters-1, 0 to Layer_3_Inputs-1) :=
  (
    (11, 4, 12, 5, 12, -11, 4, 14, -44, 6, 8, 5, 21, 1, -4, 27, 12, 26, 24, 19, -62, -21, -2, 38, 24, 3, 19, 17, 1, 29, 21, 15, -24, 5, 4, 46, 27, 3, 13, 53, 44, 17, 20, 32, -51, -12, 18, 38, 37, 26, 0, 43, 38, 54, 51, 34, -71, 0, -5, 68, 29, 27, 8, 11, 3, 40, 39, -9, -31, 26, 11, 45, 24, -10, -16, 27, 21, 27, 14, 31, -28, -4, 14, 23, 28, 5, -3, 30, 21, 36, 28, 10, -23, 12, 17, 20, 23, 29, -4, 17, -5, -5, 10, -23, -12, 20, -4, -32, -10),
    (-7, -77, 17, -19, -10, -2, -29, 13, 17, -26, -24, -25, 18, -66, -12, -22, 42, 28, -9, 48, 1, 5, -24, 8, 9, -44, -5, -32, 19, 6, -9, 23, -6, -33, -2, 26, -23, -56, 29, -28, 3, -41, -25, 6, 13, -2, 24, -1, 10, -95, 11, -26, 3, -7, -4, 17, 13, -3, -4, 43, 26, -48, -24, -27, 28, -26, -1, 11, -7, 0, -11, 27, 6, -34, 4, -21, 12, 0, -18, 14, 7, 39, 45, -3, -6, -52, 33, 8, 24, -16, -31, 28, 5, 12, 6, 11, 14, -52, 11, -2, -12, -43, -10, 27, -26, -7, -12, 31, 1),
    (4, -24, -27, -37, -20, 23, 3, 13, 2, 5, 4, 38, 14, -55, -11, 1, 4, 33, -16, -10, 20, -17, 15, -4, 6, -12, 9, -4, 3, 4, -10, 0, 24, -2, 8, -13, -36, -44, 8, -29, -13, -16, 31, -13, -4, -28, -29, 20, 10, -43, -19, 9, 9, -14, -27, -2, 22, 7, 5, -43, 12, -22, 13, -15, 3, -15, -46, -15, 36, -17, 31, -55, -44, -31, -23, 21, 21, -7, -10, -4, -4, -19, -32, 8, -17, -46, -28, -43, 14, -66, -66, -7, 28, 25, 4, -28, -1, -24, 4, -2, 5, -57, -44, 7, 20, 37, 29, -26, 2),
    (5, -59, -9, 0, -1, 35, -2, -28, 12, -1, 5, -3, -1, -25, 29, -24, -12, 11, -27, -57, -11, 6, 1, -47, 17, 4, 1, 6, -4, -11, -20, -25, 8, -4, 31, -58, -5, -51, 25, -36, -3, -44, -35, -19, -5, 20, 20, 23, -8, -51, 30, -21, -16, -33, -57, -39, -12, 41, -2, 24, 3, -14, 11, 2, -1, -1, -58, -19, -5, 29, 35, 5, -17, -32, -7, 1, -12, -8, -7, -9, -24, 13, 10, 25, -7, -31, 23, 10, -5, -5, 17, -6, -20, 8, 12, 33, 20, 5, 38, -37, 20, 1, 18, -9, 6, 13, 16, 13, 5),
    (-27, 46, -47, -18, -36, -50, 2, -25, 20, -20, -41, 18, -7, -14, -28, -48, -36, 2, -11, 5, 2, 4, -8, 56, 7, -2, -46, 8, -22, 23, -13, 19, -11, -35, 10, 20, -8, 23, 44, -5, -45, -8, -24, 6, 6, -8, 13, -86, -14, -6, 31, 19, -4, -12, -16, -3, -37, 21, 18, -51, -15, -65, 29, 12, -9, -6, -4, 26, -43, 12, -3, 21, 0, 34, 27, -7, -4, 14, -5, -12, -4, 3, 11, -28, 18, 21, 19, -1, 8, 24, -8, -1, -30, 6, -5, -23, 39, -21, -2, 11, 27, 23, -2, 2, -24, 28, 3, 32, -6),
    (0, -28, 31, -57, 15, -38, -7, 16, -17, 32, 28, 33, -6, -37, 23, 13, -18, -18, -3, -6, -68, -6, 6, 14, -15, 11, -10, 29, -8, 27, 8, 0, -39, -42, -29, -13, 26, -45, 22, -59, 13, -9, -24, 39, 48, 33, 45, 32, -1, -60, 5, -33, -13, -21, -23, -7, -20, -19, -18, -14, -35, -17, -21, 14, -54, -6, -3, 20, -38, -13, -31, 15, 29, -31, 12, -44, 26, -10, -7, 12, 44, 38, 32, 19, -7, -34, -14, -51, 6, -36, -8, -13, -42, -10, -16, 17, -35, -30, -13, 8, -3, -5, -6, 14, 9, -31, -18, 3, 11),
    (-5, -29, 4, 15, -4, 37, 16, -18, 5, 11, -37, 7, -26, -3, -1, -25, -26, -40, 16, -32, -45, -11, -31, -27, -18, -1, -33, -4, -24, 15, 6, 12, -14, -2, -5, -27, -5, -28, -16, 11, -43, -15, -2, -6, 6, -35, 6, -6, 19, -17, 14, -7, 12, -17, -19, -21, 7, 8, -6, -24, -12, -21, -41, -6, -45, 17, 8, -33, -22, 8, -34, 10, -22, -2, -43, -5, -31, -32, -11, -7, -39, -19, -63, 21, -11, -3, -28, 18, -9, 13, -32, -31, -13, -40, -10, 25, 9, -3, -4, 4, 4, -26, -3, -26, -14, -20, -30, -19, -2),
    (-15, 31, -23, 40, -16, 26, 8, -4, -31, 4, -10, -3, -22, 5, -17, 11, -16, 5, 0, 3, -38, 5, 20, 4, -9, -13, 21, 15, 5, -31, 5, -28, -5, 34, 28, 21, -5, 36, -30, 18, -4, 10, 5, -38, -27, -4, -8, -27, 11, -4, -12, 5, 8, 4, 2, -31, -46, 11, 35, -20, 15, 5, 6, -21, 11, -30, 0, -58, -28, 33, 24, 2, 18, 28, -28, 28, -15, 14, -11, -49, -12, 20, 3, -28, 31, -2, -2, 18, -8, -19, -15, -21, -4, 50, 47, -21, 23, -14, 13, 26, 15, -28, 5, -37, 11, 37, 35, 1, -7),
    (13, 28, -5, -46, -12, 4, -12, -17, 12, 9, 43, -33, 29, 14, -38, -8, -10, -36, -17, -13, 32, 22, 36, -60, 17, 22, -11, 28, -17, -11, -20, -14, 4, -23, 13, -40, 20, 14, -34, -33, -14, -26, -37, -3, 22, 33, 43, -38, 37, 26, -38, -37, -14, -27, -41, -42, 22, 1, 49, -44, 27, 21, -7, 8, -11, -10, -5, -24, -4, -14, -5, -14, 15, 4, 1, -22, -12, -28, -13, 12, 13, 28, 42, -28, 20, 4, -5, -10, 7, -10, -12, -34, 17, 33, 31, -3, 20, 6, 0, 15, 3, 3, 18, -27, -17, -10, -8, 7, -6),
    (-20, -4, -5, 10, 11, -49, 15, -47, -23, -1, 5, 18, 24, 12, 26, 30, 12, -34, 39, -49, -70, 33, 0, 29, 43, -4, 3, -1, -20, -43, 20, -4, -28, -14, 29, 17, 6, -13, -21, -15, -48, -47, 20, 13, -36, -15, -17, 41, 29, -12, -28, 39, 4, 0, 42, 41, -58, -25, 10, 23, -15, 13, -3, 15, 31, -10, 23, 31, -86, -31, -20, -13, -44, -51, 13, 9, -5, -30, 22, 34, -33, 23, 13, -4, -12, -64, 25, 19, -66, -15, 45, 21, -31, -15, -1, 3, -32, -42, -4, 19, -6, -8, -3, 12, -33, -28, -48, -33, -6),
    (1, -45, 0, 29, -19, 27, 4, -5, 12, -20, -23, -5, -14, 12, -8, 5, -19, 7, 0, -19, 17, 19, 12, -16, -20, 47, 39, 39, 3, -8, -13, -13, 22, -3, 5, -33, -7, -1, 7, 14, 8, 17, 10, 31, -9, -51, -27, 39, -22, 40, -11, 29, 8, 25, 26, 14, -15, -15, -6, 2, -32, 43, -31, -27, 6, -46, 4, -44, -16, -20, 21, -31, 2, 3, 11, 6, -53, 10, 56, 36, -1, -12, -15, 39, -34, 31, 35, 4, -45, 19, 16, 39, -18, -7, -38, -20, -14, 9, 4, -16, -28, -19, -32, 8, -1, 22, 9, -34, 0),
    (-75, -39, -28, -21, -32, 2, 6, -19, -11, -1, -59, -55, -48, -53, 19, 0, -35, 4, 45, -17, -30, -1, -32, -26, -32, -19, 2, 3, -36, -13, 31, 16, -19, 5, -35, 34, -9, -8, 8, 45, -39, 30, -12, 12, 13, 5, -4, -37, -15, 28, 38, 35, -1, 18, -25, 42, 4, 9, -7, -20, 11, 40, 28, 16, 25, 6, -12, 18, -2, -1, -1, 3, -11, 20, 12, 0, 20, 28, 8, 4, 24, -9, -16, -11, -10, 12, 5, 27, 39, 32, 27, 26, -3, -6, 12, -5, 20, 26, -1, -5, 33, 18, 29, -3, -21, 7, 32, -20, -3),
    (-20, -6, -17, -59, -22, 14, 4, 32, 12, -9, 36, 14, -5, -1, 6, 2, 3, 19, 24, 21, 25, -5, 27, 34, 15, 13, 3, -26, 4, 14, 29, -16, 28, 35, 19, 30, -17, 0, -18, -2, -9, 13, 13, 13, -16, -25, -12, 3, -12, 12, 13, 28, -4, 44, 33, 33, -12, 2, 27, 46, -17, 10, 27, -9, 4, 28, 32, 17, 12, 18, -2, 28, -21, -19, 19, 16, 22, -18, 17, 32, -10, -15, 6, 27, -19, 11, 11, 0, 13, 5, 44, 17, -4, 23, 9, 31, -3, 18, 8, 17, 2, 5, 22, -16, 6, 5, 21, 3, -13),
    (-26, 3, -17, -31, 3, -28, -11, -25, 9, -28, -13, 8, -16, 20, -6, 13, 1, -29, 3, -7, -1, -9, 1, -5, -7, 37, -27, -15, 10, 8, -5, 13, -6, -6, -12, -39, -42, 24, -62, -11, -8, -65, 13, -6, -5, 0, -24, 24, -40, 23, -18, -15, -13, -23, 27, -10, -17, -22, -30, 6, -33, 19, -31, 5, -36, -3, 1, 4, 14, 11, -10, -23, -17, 4, 19, 35, -60, -3, -13, -6, 16, 1, -5, -39, -13, 9, 26, 17, -47, -11, -12, -15, 4, 38, 23, -76, -10, -21, 40, 14, -5, -16, 3, -12, 22, 38, 39, -40, -9),
    (-9, 27, 4, -22, 23, 51, 28, 31, -31, -21, -6, 9, -12, 8, -17, 6, 23, 42, 19, 80, 11, -36, -4, -1, -21, 16, 12, -18, 23, 20, 7, 47, 12, -20, 8, -15, -12, -12, -12, 18, 30, 14, 50, 22, -21, -3, -48, -11, -22, -36, 0, 16, -19, 37, 30, 17, 2, -3, 1, -63, -23, -56, -4, -18, -12, 10, -5, 10, -12, 17, -29, -25, -2, -12, -1, 29, -4, 20, -15, 24, 12, 28, 36, -15, 9, -24, 20, 26, -9, 1, -13, 26, 41, 4, 35, 13, 19, -10, 20, 28, -13, -7, -27, 29, 21, 18, 2, 22, -6),
    (7, 31, 18, 57, -32, 0, 5, 10, 6, 14, 41, -4, 6, 20, 4, 51, -20, 12, -5, 1, 2, -6, 25, -5, 14, 5, 4, 2, 4, 16, -2, -11, 4, 13, 20, -2, 4, 34, 24, 54, -31, 53, 16, -12, -40, 19, 10, 29, -5, 17, 8, 54, 11, 27, 26, -22, -73, 1, -12, 37, -1, 18, 4, 17, 6, -5, 9, 1, -44, -22, -26, 23, -21, 13, -6, 40, -24, 7, 34, 8, -56, -7, -44, 34, -30, 20, -8, 29, -13, 55, 33, 38, -100, -31, -35, 27, -30, 28, 17, 11, -17, 41, 17, 49, -100, -43, -37, -19, 7)
  );
  ----------------
  CONSTANT Layer_4_Columns    : NATURAL := 16;
  CONSTANT Layer_4_Rows       : NATURAL := 16;
  CONSTANT Layer_4_Strides    : NATURAL := 2;
  CONSTANT Layer_4_Activation : Activation_T := relu;
  CONSTANT Layer_4_Padding    : Padding_T := same;
  CONSTANT Layer_4_Values     : NATURAL := 16;
  CONSTANT Layer_4_Filter_X   : NATURAL := 3;
  CONSTANT Layer_4_Filter_Y   : NATURAL := 3;
  CONSTANT Layer_4_Filters    : NATURAL := 24;
  CONSTANT Layer_4_Inputs     : NATURAL := 145;
  CONSTANT Layer_4_Out_Offset : INTEGER := 6;
  CONSTANT Layer_4_Offset     : INTEGER := 0;
  CONSTANT Layer_4 : CNN_Weights_T(0 to Layer_4_Filters-1, 0 to Layer_4_Inputs-1) :=
  (
    (12, 4, 18, 1, 9, 17, 2, 4, 4, 26, -2, -12, 6, -2, -16, 12, 41, -11, -5, 11, 20, 15, 1, -3, -12, 53, 21, -4, 12, -11, 9, -5, -18, -8, 32, 8, -39, 25, -18, -21, -8, 1, 4, -24, -28, -35, 17, -24, 21, 9, -9, -1, 34, 12, 21, 15, -9, 19, 27, 5, 20, 16, 15, -1, 44, -10, -15, -4, -18, 23, 31, 3, -28, 25, 18, -29, 12, -4, 20, -9, -44, 9, -3, 4, -36, 20, 24, -8, 4, -10, -37, -31, -27, -46, -1, -25, 20, -1, -35, -8, 28, 12, 4, -1, -14, 30, 39, 20, 17, 16, 18, 15, -16, -12, -14, -18, -21, -8, 13, -16, 3, 19, 4, 3, -40, -6, 22, 3, -62, -11, -11, -35, -43, 24, 17, 24, 28, 4, 6, -43, -20, -55, -29, -2, -3),
    (-36, 25, 16, 2, -45, 20, 1, -1, -38, -26, -27, -23, 4, -10, -8, -59, -19, 24, 30, 28, -29, 26, -31, -30, -38, -39, -35, -11, -34, -36, 12, -22, -30, 22, 10, 14, -22, 23, -4, 4, -5, -5, 5, -23, -33, -33, 13, -14, -22, 33, 0, 40, -28, 28, -16, -3, 3, -31, -14, -8, 19, -26, -6, -7, -42, 40, 28, 48, -32, 36, 7, 7, -4, -33, -17, -13, 23, -20, 22, -1, -29, 27, 3, 7, -22, 4, 11, -2, -7, -8, -35, -21, 4, -10, 24, 0, 11, 38, 12, 13, -1, 26, -25, -5, 8, 54, -16, -1, -2, -20, -3, 24, 5, 35, -3, 25, 1, 7, 17, -9, 4, 28, -2, 11, 4, -7, 21, 0, -1, 6, -14, 6, 11, -11, 2, 14, -7, -2, 7, 6, 4, 27, 8, -5, 6),
    (17, -3, -5, 34, 36, -6, -28, 17, 8, 25, -13, 17, 17, 16, 11, 27, 28, -4, -4, 33, 29, -24, -6, 35, -8, 42, -11, -3, 0, 20, 20, 22, 28, -12, 1, 24, 4, -8, 19, 14, -11, 22, -13, -21, 22, -5, 34, -4, -4, -18, -8, 12, 10, 25, -7, 16, -15, -15, -10, 4, 12, 3, -3, 13, 15, -24, -20, 31, 21, 12, 12, 16, -8, 40, -5, 12, 9, 24, 29, -5, 17, 0, -7, 25, 14, 13, 53, 34, -5, 33, -18, 4, 3, 2, 1, -36, 4, 11, 10, 8, 0, 26, 50, 3, 5, 4, -18, -32, 9, -15, 4, -15, 10, 12, -16, -11, 22, 9, 31, -2, -25, 13, 13, 1, -3, -4, -2, -27, -20, 27, -10, -12, -4, 5, 37, 0, -27, -12, 13, 28, 16, 10, -16, -19, -23),
    (-6, -6, 12, 13, 0, 40, -54, 19, 28, -17, -4, -10, 20, 12, -11, -3, -25, -21, 42, 14, -29, 25, 0, 4, 3, 23, -13, -21, -14, -9, 7, 6, -16, -11, 12, -11, 4, -29, 30, -3, -1, 16, -32, 1, -32, -19, -13, -8, -24, -6, 23, 4, -14, 26, -19, 34, 30, -26, -12, -30, -14, -40, -11, -8, -23, -25, 12, -13, -68, 15, 1, -21, 12, -43, -31, -14, -23, -18, -47, -10, 48, -27, -4, -16, -33, -18, -27, -9, -24, 14, -16, 46, -13, -20, 9, 9, -27, 2, 25, 16, -12, 25, 6, -10, 28, -20, -29, -34, -8, -57, -16, -29, -1, -30, -9, 7, -48, 13, 13, -46, -7, -3, -4, -2, -6, -33, -16, 3, 35, 2, -13, -13, -18, -10, -22, -23, -39, -9, 23, 29, 29, -11, 21, -5, 14),
    (16, -11, -13, -3, 1, 0, 11, -1, 15, -17, -42, -9, -9, -10, -21, 1, -1, -15, -17, 1, -5, -22, 43, -16, 12, -11, -23, -23, 1, -20, -33, -4, -16, -25, 10, -17, -23, -33, 18, -5, 12, -10, 16, -4, -8, -15, -10, -11, 34, -40, -4, 2, 4, 36, -3, 33, 16, -20, -49, -24, 9, -21, -37, -11, 48, -30, -21, 13, 4, -6, 42, 28, 19, -6, -52, -53, 17, -50, -52, 3, 38, -28, -2, 0, -9, -34, 15, 4, 12, 15, -13, -29, 4, -12, -12, 12, 21, -19, -18, -9, -17, 11, -8, 13, -11, -12, -5, -10, -1, -18, -8, -13, 37, -21, -15, -2, -15, 11, 2, 53, 24, -16, -21, -38, 30, -10, -28, -14, 23, -33, 4, 1, -6, -4, 10, 23, 31, 1, -4, -21, 13, 14, -13, -22, -10),
    (-4, -2, -9, 6, -38, -5, -1, -23, -20, -4, -10, -18, 9, -28, 5, -18, -38, 9, 1, -21, -29, -4, 6, -33, -3, 10, 7, -12, 2, -14, -14, -38, -18, -8, -7, -9, 3, -5, 26, -18, -2, -11, -21, 11, -2, 7, -18, 2, -21, 1, -6, 5, -19, 6, -3, -15, -2, 10, 26, -32, -2, -16, 16, -14, -48, -20, 15, 12, -21, 5, -10, -15, 12, -14, -8, -32, -11, -11, -4, -3, -30, -46, 20, -7, 7, 9, -12, 25, 25, -9, 1, 9, -13, 12, -20, 4, -10, -8, 20, 30, -8, -21, 4, 4, 24, -36, 2, 15, 4, 17, 16, 14, -13, -34, 65, 42, -10, -1, -23, 12, 42, -61, -27, -20, 19, 12, -4, 45, -6, -45, 46, 23, -4, 4, -16, 2, 22, -28, -10, -12, 13, 15, 2, 36, 6),
    (9, -10, -14, 2, -22, -19, 9, -21, -45, 32, -5, -57, -5, 4, 9, 2, 30, -42, -26, 37, 3, -19, 55, -16, 4, 50, -19, -30, -3, -5, 17, 14, 19, -38, -17, 32, -8, -56, 19, 3, 9, 28, -6, 19, 20, -18, 29, 33, -39, 13, 2, -15, 3, -21, 51, -19, -31, 63, 31, -31, -6, 6, 9, -13, -16, 14, 4, 14, 5, 4, 26, 0, -26, 24, -9, -32, -21, 6, -4, 11, -15, 12, -4, -32, 27, -2, 31, -7, -33, 4, -17, -19, -59, -2, 10, -10, 21, 3, -14, 21, 30, -12, -2, 28, -9, 44, 6, 22, 2, 19, 15, 25, 21, 5, -7, 33, 22, -2, 16, 14, -16, 36, 14, 8, 8, 28, 0, 10, 0, 10, -2, 13, 13, -18, -10, -13, -26, -8, 18, -15, -25, -11, 23, -23, 4),
    (-3, -39, 8, -20, 10, -11, 8, -8, -4, 9, -6, 5, 17, -6, 4, 2, -12, -14, 9, 21, 25, 83, -7, 9, 2, 5, -17, -25, 3, 16, -12, -27, 12, -8, 29, 28, -27, 54, -33, 39, 36, -35, -20, -36, 12, -21, -34, 3, -23, -39, -9, 9, -10, -8, 28, 6, -18, 14, -25, -31, -24, -14, -20, -15, -10, -27, 24, 29, -44, 42, -7, -4, 17, 8, -39, -65, -13, -43, -41, -15, -12, -6, 21, 8, -47, 37, 2, -10, 13, 4, -19, -43, 16, -45, -21, 1, -24, -27, 7, 1, -16, -7, 29, 0, -14, 1, -13, -46, -28, -59, -46, -22, 6, 9, 12, 15, -21, 20, 17, -17, -30, -5, -33, -65, -15, -60, -52, -3, 10, -4, 9, 21, -22, 11, 2, 5, -12, 4, -6, -37, 20, -11, 8, 11, 11),
    (-5, -36, 43, 45, -37, 47, -19, 9, 28, -31, -33, -11, 6, -32, -18, 21, -6, -5, 62, -2, -24, 13, 18, -13, 9, 13, -18, -10, 8, -12, -22, 23, 10, 7, -18, 0, -14, 6, -12, -69, -4, 10, -26, -21, -18, -36, 12, 4, -4, -15, 31, 13, -35, 27, 26, -35, -12, -13, -10, -10, -13, -42, -40, -4, 19, -33, 44, 1, -4, 38, 5, -48, -26, 26, 12, -26, 29, -24, 8, -11, -10, 5, -11, -4, -13, 12, 4, -60, -33, 5, 19, -29, -42, 0, -12, 2, 21, -29, -25, 0, 3, -12, 44, -21, -19, 36, 3, -5, 4, 10, -5, -16, 25, -16, -14, 28, 3, -12, 21, -24, -37, 21, 19, -21, 5, 15, 32, 3, -25, 5, -6, 14, -21, -38, 26, 3, -18, 20, 2, -21, -17, 31, 17, 10, 28),
    (-16, 10, -2, -16, -19, 8, -10, -25, -19, -6, -15, -17, 4, -20, -10, -9, 11, 22, 8, 34, 0, -65, -42, 5, 21, -8, 22, 4, 34, -1, 11, 15, 11, 4, 6, 9, 13, -23, -37, 25, 8, -4, 52, 6, 17, -4, 27, 22, -5, 28, -13, -20, 4, 8, 20, -2, -59, -3, -1, -35, -1, -14, -16, -46, 38, 38, -14, -4, 9, -25, 3, -11, -27, 4, 34, 20, 2, 3, 12, 0, 9, 12, -1, -7, 38, 0, 7, -3, 10, 19, 44, 16, 13, 28, 21, 12, 0, 20, -25, -24, 6, -11, 6, -22, -53, -23, 21, -6, 0, 3, -13, -28, 20, -9, -19, 4, 21, 7, -6, -13, -9, -12, 21, 12, 23, 21, 13, -9, -4, -9, 6, -14, 20, 3, 41, -4, 12, -16, 13, -12, -5, 15, -2, -3, -11),
    (-21, -6, -7, -19, -13, -4, 33, -8, -15, -20, -4, -18, -19, -12, -6, -72, -35, -13, 26, -16, -3, -51, 27, 25, 26, 0, -12, 1, -17, 11, -40, -24, -6, 1, 1, -12, 3, -51, 35, 5, 14, 24, -4, 5, 12, 10, -16, -18, -16, -3, 36, 48, -10, -21, 51, 12, 21, 20, -38, -37, 5, -1, -32, 11, 20, -28, 66, 36, 13, -44, 40, 6, 28, 28, -33, -24, 4, 11, -31, 50, 27, -1, 2, -4, 4, -24, -17, 9, 4, 1, 3, 10, 7, 9, 14, 18, 1, -6, 39, 16, 3, 15, 8, 23, 2, 16, -33, -19, -8, 6, -41, -15, 43, -24, 35, 19, -5, 13, 2, -13, 12, 31, -29, -3, -8, -29, 6, 12, 28, -12, -62, 6, -18, -9, 23, -28, -17, 8, -6, -1, -15, -12, 11, 12, -10),
    (4, -40, -12, -7, -18, -25, -7, 11, -7, -22, 12, 18, 5, 2, 15, -25, -13, -24, 13, 24, -4, 30, -35, 22, 28, -67, -16, 18, 13, 4, -1, 4, -27, -27, -16, 12, -34, -25, -33, -10, 20, 2, -2, -14, -14, -2, 11, 31, -18, -42, 1, 12, -37, -30, -3, 1, 0, -1, 10, 6, 4, -13, 22, 6, -66, -11, 52, 22, -50, 36, -29, 0, 8, -77, -2, -16, 12, -55, -29, 0, -26, -19, -29, -11, -58, 21, -17, -49, -10, -15, -24, 4, -36, -12, -50, 21, -7, -29, -3, 18, -12, -38, 24, 16, -3, 13, -8, -7, 20, -22, 3, 3, -28, -47, 16, 23, -30, 9, -16, -31, 21, -5, -11, -38, -12, -56, -60, -22, 33, -55, -106, -21, -24, 23, 24, -26, -21, -4, -22, -11, -34, -82, -52, 14, 38),
    (-21, -26, 2, -7, 11, -18, -42, 14, 26, -41, -4, 13, -8, 3, 5, 3, -17, -60, 38, -1, -5, -42, -49, 13, 49, -46, -13, 5, -4, -2, -6, 20, -4, -41, -20, -22, 3, -50, -1, 3, 11, 11, -1, 19, -12, 18, -3, 26, -30, -37, 20, 10, 6, -1, -15, 22, 28, -43, -35, 12, -1, 14, -24, 29, -13, -64, 47, 13, -21, -28, -46, -9, 32, 9, -29, 6, -13, 2, -30, 45, 3, -44, -28, -8, -10, -45, -1, -12, 22, 16, 14, 5, -20, 3, 1, 21, 6, -5, -2, 14, 13, 22, 11, -10, 19, -4, -21, -12, 4, -28, -41, 15, 28, -13, -9, 43, -19, -24, 26, -10, -9, 43, -7, -20, 5, -10, 5, 12, 22, -2, -66, 4, -10, -44, 8, 2, -27, 19, 12, -23, 7, -13, 14, -17, 6),
    (-2, -22, 24, 5, -37, -3, 29, 5, -62, -21, -13, -27, -12, -4, -50, -43, -38, -2, -14, 23, -5, 0, 41, 11, -5, 8, 22, -23, 11, -5, -20, -1, 2, 15, -34, -5, -7, -25, -46, 2, -28, -5, 26, 20, -19, 16, 6, 11, 3, -34, -28, -12, 31, -83, 50, -37, -22, 7, 7, -28, -5, 30, -4, -33, -21, 8, -33, -5, 12, -41, 32, -24, -40, 52, 43, -4, -17, 13, 14, -10, -12, 10, -29, 6, 4, -5, 11, 20, -47, 13, 54, 7, 6, 29, 30, -5, 9, -24, -7, -10, 26, -67, -1, 14, -12, -5, 30, 19, -1, 40, 28, -9, 11, -18, 4, -4, 25, -14, -26, 21, -1, -15, 8, 20, -20, 48, 20, -3, 5, -5, 8, 21, 20, 19, -11, 37, 4, 18, 21, 27, 15, 36, 21, 12, 12),
    (-44, 33, 21, -2, 10, -11, -16, 11, 23, -4, 43, 6, -20, 21, -5, -30, -37, 32, 14, 9, 19, -19, 1, 11, 36, -18, 34, 16, 7, 37, 4, -21, -12, 21, 8, 10, -6, -8, 19, 9, 16, -26, 12, 7, 3, 12, 2, -54, -6, -4, 19, 20, 50, -31, -46, -11, 24, 10, -5, 24, 3, 62, 24, 34, 4, 14, -9, 13, 70, -57, -31, -4, 7, 13, 23, 39, 9, 46, 51, 29, -13, -4, -29, -5, 18, -29, -28, -4, 3, 12, 21, 22, 28, 26, 16, -5, -4, -17, -10, -13, 38, -13, -13, -6, 5, 4, 14, 28, 9, 23, 18, 12, -3, 13, -35, -48, 41, -30, 1, -15, -30, 30, 22, 44, 5, 29, 15, -4, -21, 9, 5, -46, 8, -13, -9, -15, 4, 16, 10, 2, 11, 22, -11, -37, 5),
    (2, 56, -22, -28, -27, 8, -17, -7, -50, -7, 11, 8, -3, -20, -4, -29, 11, 32, -13, -8, -29, 64, -19, -6, -21, -50, -32, -39, 3, -47, -24, -26, 12, 32, -3, 9, -6, 8, -25, -4, -4, -23, -21, -18, 32, -16, -23, -7, 2, 35, -25, -13, 1, 4, -14, -35, -45, -9, -14, -10, 21, -12, 10, -35, 28, 39, -12, 0, -50, 53, -12, 11, -52, -3, -28, -47, 27, -68, -32, -14, 27, 10, -6, 11, -44, 20, -5, -4, -26, -21, -27, -25, 44, -40, -20, 14, -4, -2, 29, 9, -11, -16, -22, -8, -23, -7, -5, -13, 25, -14, 2, -15, 20, 15, -2, -3, -19, 2, 28, -10, -34, -10, -12, -15, -6, -33, -12, -4, 29, -2, 1, 11, -30, 37, 1, 30, 7, 2, -23, -14, 15, -47, -22, -7, 24),
    (-53, 16, 7, -24, -1, -56, 66, 2, -54, 19, 4, -5, -38, 24, -4, -13, -30, 40, 10, -24, 25, -29, 19, -8, -39, 13, -9, 4, -24, -18, 4, -17, 11, 27, 12, -18, 18, -28, -16, -18, -44, 14, 8, 6, -12, -11, 3, 7, 12, -10, -10, -5, 27, -46, -2, -2, -29, 25, -8, 24, -20, 1, 10, 9, 37, 21, -1, -8, 49, -33, 4, 17, -48, 8, 4, 25, -3, 18, -12, -12, 46, 7, -21, -2, 28, -16, -33, 14, -19, -6, 23, 24, 11, 12, -1, -12, 14, -7, 16, -9, -20, -3, 2, 20, 12, -1, -37, -13, 12, -50, -24, -10, 26, -4, 7, 13, 2, -5, -11, -10, 16, -15, -24, 2, 13, -25, -12, 4, 21, -4, -7, 7, 3, -10, -35, -13, 3, -12, -4, 0, 24, 10, 1, 7, 1),
    (22, 14, 10, -2, 18, 28, -14, 31, 8, 20, -10, -4, -12, 12, -17, -8, 30, 20, 13, 13, 11, 28, 25, -5, 3, 4, -24, -21, -14, -12, -13, -20, 11, 18, -38, -32, -24, 8, 9, -31, -5, 49, -19, -12, -26, -57, 4, 7, 4, 40, -1, -13, 33, 36, -34, 30, 18, 19, 3, -4, -9, 36, -17, -22, 8, 44, 7, -12, 52, 43, 14, 40, 7, 4, -5, -5, 20, 28, -22, -19, -4, 18, -34, -3, -7, -6, 39, 4, 12, 15, -55, -38, 9, -43, -27, -13, -10, -5, 6, -24, 21, 7, -25, 21, 4, -10, -2, 11, -13, 25, -11, -31, 4, 0, -7, -12, 37, 13, -19, 33, 16, 1, 5, 4, -9, 19, -12, -28, 4, 18, -30, -4, -3, -31, -17, -15, 18, 11, -33, -13, -35, -40, -7, 4, -10),
    (-33, -5, -31, -34, -13, 13, -60, -18, 13, -15, 16, -10, -4, 7, 9, 4, -20, 17, -14, -19, -25, 40, 1, -13, 12, -7, 34, 9, -10, -9, -3, -8, -25, 0, -1, -10, -15, 37, -1, 0, -4, -13, 32, -8, 22, 13, 4, -8, -21, -28, -10, -6, 7, 15, -28, 19, 17, -7, 17, 13, -10, 6, 2, 3, -35, -24, 12, 18, 7, -2, -17, 10, 39, -20, 19, -7, -9, 6, -1, 3, -12, -16, 45, 26, 3, 4, -24, 13, 39, 9, 15, 0, 21, 22, 1, 44, 4, -26, 6, 8, -3, 7, 14, 0, 6, 9, -6, 0, 18, 20, -1, 23, -28, 0, 14, 9, 7, 7, -12, -2, 36, 4, -24, 6, 8, 12, -19, 27, -8, -3, 19, 21, -11, 8, 13, 15, 27, 15, -17, -14, 13, 23, -14, 16, -16),
    (3, 20, -28, -26, 5, -20, 35, -39, -43, 1, 8, -8, 2, -20, -10, -13, 28, 35, -35, -22, 19, -17, -17, -17, -48, -6, 10, 18, -12, 18, -14, -7, 24, 34, -31, -12, -3, -19, 5, 8, -21, -14, -3, -4, 34, 8, -13, -20, -34, -5, 16, -10, -5, -13, -1, -31, -35, 43, -6, -20, 5, -29, -37, -14, 31, 44, -38, -12, 37, 3, -11, -19, -28, -13, 44, 20, 26, -8, 16, 7, 9, 25, -17, -24, 24, 10, -13, 4, -6, -35, 11, 12, 40, 13, -6, -1, -33, -3, 7, 9, -1, 3, -4, -13, -38, 10, -20, -5, -4, -6, -30, -20, 30, 47, -19, -5, 15, -1, -17, 23, -33, 8, 41, 12, 11, -10, 21, -6, 3, 16, -4, 2, 0, 4, -4, 27, -3, -11, 27, 10, 12, 14, 9, -12, 4),
    (22, -10, -26, -21, 12, -43, -1, -9, 12, -3, -4, 2, 12, -2, 19, -4, 24, -3, -29, -35, 7, -5, 3, 8, 6, -6, -5, -10, 31, -4, -12, -42, 4, 10, -11, -4, 8, 10, 0, 8, 0, -11, -6, -16, 20, -3, -20, -27, 28, 19, -35, -39, 19, -28, -2, 20, 7, -20, 25, -4, 9, -11, -3, -14, 30, 9, -35, -50, -4, -13, 2, 32, 24, -28, 18, -12, 23, -4, -13, -62, 12, 17, -28, -20, 1, 7, -1, -1, 7, -24, 20, -3, 16, -11, 9, -50, 26, 7, -6, -2, -2, -13, -39, 29, 16, -1, 12, 3, 21, 8, 5, -22, 24, -10, 5, -20, -9, -12, -23, 23, 18, -28, 27, 8, 20, 9, 7, -52, 2, -4, 10, -6, -5, -6, -39, 1, -4, -41, 7, 9, 28, 3, 3, -24, -16),
    (25, -15, 5, 18, 6, -19, -13, 12, 12, 5, -9, 12, 7, 20, 20, 42, 16, -38, -1, 11, 4, -41, -15, -11, -3, 19, -1, -2, 9, -1, 15, 19, 20, -35, -19, 7, 6, -42, -4, -25, 4, 14, 10, -10, -1, 4, 8, 8, 52, -4, -12, 1, 21, 3, 14, -3, -17, 46, -4, -14, -13, -14, 18, 32, 34, -7, 27, 16, 0, 4, 9, -5, -35, 47, 4, -7, -1, -31, 34, 17, 17, -10, -6, -13, -1, -29, 28, -29, -34, 29, 24, 19, -22, -15, 23, 20, 15, 15, -50, -28, 7, 6, 39, 8, -19, 21, -7, -8, -30, -28, 4, -30, -3, 32, -41, -2, 6, 50, 23, -2, -14, 36, -17, -18, -26, -20, -21, -45, 4, 28, -23, 4, -19, 35, 39, -24, -28, 25, -34, 8, -68, -45, 11, -28, 1),
    (10, -10, -22, 10, -12, 8, 16, 30, 13, 10, -28, -21, 16, -26, -24, -30, 28, 8, -13, 11, 31, 2, 12, 7, 21, 30, -44, -2, 8, 7, -14, -4, 19, -9, -13, 9, 14, -4, -21, 8, 9, 1, -14, -10, 20, 12, -18, 6, -36, 12, -1, -20, -8, -14, 13, -30, -4, 2, 4, -26, -11, 3, -23, -49, 12, -3, -33, 17, -24, 0, 3, 3, 5, 20, -37, -25, -6, -27, -30, -4, 40, -41, -43, 27, -12, -5, -13, 23, -4, 11, -41, -4, 28, -28, -20, 7, -57, 16, 28, 13, -10, -11, 6, -32, 11, -14, 29, 1, 18, 24, -9, -4, -53, -6, 20, -21, -25, 1, 12, -44, 6, -36, 5, -7, -16, 20, -19, -3, -29, 13, 4, -37, -11, 3, -9, -15, 1, -25, -11, -13, -29, -37, -45, 1, -8),
    (-21, 30, 6, 12, 14, 3, 29, 2, -38, 28, 19, 3, -5, 24, 2, -30, -22, 47, 31, 10, 31, -23, 14, -12, -28, -12, 12, 5, -42, 6, -1, -15, -13, 21, 15, -1, 25, -9, 1, -37, -31, -4, -2, -13, -43, 14, -17, -10, 24, 18, 4, 4, 27, 40, 22, 30, -25, 48, -20, 25, -12, 30, -4, -22, 23, 14, -6, 21, 19, 38, 22, 28, -10, 23, -3, 20, -32, 15, -4, -60, 4, 5, -10, -4, 22, -6, -7, 1, 11, 15, -2, 0, -29, -17, 5, -47, 12, 33, 10, -5, 1, 28, 16, -4, 16, 1, -12, 4, -23, -4, -10, -19, 6, 61, 2, -12, -18, 42, 21, 23, 9, 4, -28, 4, -11, -38, -29, -47, 24, 6, -6, 11, -44, 22, 6, 11, -10, -32, -30, -34, -24, -48, -35, -45, 1)
  );
  ----------------
  CONSTANT Layer_5_Columns    : NATURAL := 8;
  CONSTANT Layer_5_Rows       : NATURAL := 8;
  CONSTANT Layer_5_Strides    : NATURAL := 2;
  CONSTANT Layer_5_Activation : Activation_T := relu;
  CONSTANT Layer_5_Padding    : Padding_T := same;
  CONSTANT Layer_5_Values     : NATURAL := 24;
  CONSTANT Layer_5_Filter_X   : NATURAL := 3;
  CONSTANT Layer_5_Filter_Y   : NATURAL := 3;
  CONSTANT Layer_5_Filters    : NATURAL := 32;
  CONSTANT Layer_5_Inputs     : NATURAL := 217;
  CONSTANT Layer_5_Out_Offset : INTEGER := 6;
  CONSTANT Layer_5_Offset     : INTEGER := 0;
  CONSTANT Layer_5 : CNN_Weights_T(0 to Layer_5_Filters-1, 0 to Layer_5_Inputs-1) :=
  (
    (6, -9, -20, -39, 5, -3, 9, -35, -23, 6, -11, 29, -28, 20, 14, 4, 21, -3, -10, 37, -5, -12, -12, -27, 12, -32, 16, 50, 12, -8, -39, -6, 2, -3, 3, 20, 17, 12, -24, -5, 11, 31, 5, 44, 17, -13, -30, -43, 21, -20, -5, 19, 4, -4, -5, -4, 16, -4, 13, 4, 22, -35, -12, 4, 3, 4, -11, 1, 3, 20, 0, -42, -12, -21, -16, -14, 4, -4, -10, -20, -9, 5, -10, -4, -29, 15, -6, -7, 20, 25, 21, 3, 2, -22, -2, -16, 22, -40, 19, 21, 23, -19, -45, 5, 28, 4, 19, -20, -3, 8, -29, -20, 18, 46, 13, 10, 4, -12, -20, -49, 15, -3, 12, -12, 7, -8, -37, 5, 24, -29, 6, -6, 26, -35, -13, -47, -12, 17, -22, 5, 1, 1, 14, -36, -9, 13, 19, -14, 12, -22, -13, -4, 3, 10, 8, -7, -2, 5, -17, -6, -3, 19, 12, -11, 11, -21, 20, -7, 18, 7, 17, -3, 19, -5, -35, 2, -11, 19, 19, -15, -4, 0, -2, -8, -2, 22, 20, 4, 14, -15, 11, -21, 11, 4, 5, 9, -20, -3, -21, 19, -5, -32, 19, 12, -5, -14, -12, -54, -4, 17, -2, -18, 0, 3, 2, -32, -13),
    (12, -13, 13, -31, 25, 25, 20, 24, -3, -11, 18, -13, 7, -46, -2, 0, -44, 5, 14, -43, -14, 10, 25, 16, 7, 12, 13, -46, 19, 36, 20, 21, -19, -10, 23, -35, 12, -23, 4, -4, -12, -4, 21, -53, 3, 13, 12, 1, 2, 3, 8, -21, 19, 34, 7, 7, -16, -10, 23, -28, 7, 9, 7, -12, 5, -14, 14, -14, -3, 11, -4, 7, -26, 2, -15, -27, 3, 3, 13, 15, -11, -1, 0, -6, -44, -12, -18, 11, -31, -15, -21, -21, -15, -12, 18, 22, -15, 0, -16, -37, 18, -1, 31, 4, 4, -9, 6, -4, -17, -16, -11, 33, -29, -13, -5, -38, -28, 7, 12, 11, -7, 16, -24, -26, -7, 17, 28, -11, 4, -20, 31, -25, 5, -37, -5, 26, -9, -23, -27, -14, -19, 13, 0, 25, 5, 1, 4, 34, 12, -14, -9, -10, 23, -16, -5, 15, -17, -31, -29, 20, -3, 38, -34, 16, -1, -5, 2, 27, -20, -2, 4, -16, 5, -27, -15, -27, 11, -18, -24, -13, -25, -28, -31, 3, -35, 1, -17, 16, -8, -4, 23, -16, -2, -2, -14, -18, -8, -14, 2, -11, 31, -3, -14, 9, -11, 9, -5, 10, -12, -2, -25, 2, 2, 9, 36, -29, -6),
    (28, 13, 11, -11, 2, 15, -13, 37, 2, 16, 30, -20, -6, -4, 12, -25, -47, 32, -7, -38, -28, -2, 11, 7, 37, 9, -4, -17, 3, 28, 14, 8, 3, -10, -23, -2, -4, 18, -25, -2, 32, -7, -20, -15, -31, 35, 25, 9, 11, -19, -43, -14, 7, -3, 20, -12, -22, -14, 13, -17, -27, 9, 0, -14, 37, -20, -16, 12, 8, -7, -16, 3, 13, 22, -22, -20, -10, 16, 25, 21, -6, -3, 10, -20, -36, 5, -6, -21, 5, 13, -34, -15, -16, 8, 20, 11, 10, -25, -11, 4, 21, -1, -8, -12, -16, -17, -4, 25, -47, 29, -27, 41, 27, 7, -6, 8, -19, 20, -1, 17, 24, -42, -20, 18, 32, 4, 5, 12, -11, 8, 20, 7, 17, 2, -23, 23, 34, 7, 13, 40, 8, -34, -24, -18, -18, 12, -18, -8, -38, 0, 23, -2, 5, -14, -1, -20, -14, -3, -22, 18, 20, -22, -5, 2, 7, -4, 13, 8, 17, -13, 2, -7, 38, 11, -3, -25, -13, -4, 4, 6, -33, 28, -26, 35, 14, -2, -3, 28, -4, -10, -12, -10, 17, -23, -5, 22, 27, 11, -16, -4, 28, -1, 0, -5, 6, -3, -14, 14, -6, -2, -13, 3, -6, 2, -37, -7, -1),
    (13, -7, 20, -12, 6, -11, 4, 6, 12, 1, -11, -4, 7, 18, -3, -8, 13, 4, 1, 5, 4, -29, 37, -4, 8, -8, 3, -6, 15, -15, -3, -11, -3, -4, 2, -8, 4, 29, 3, -9, -6, 8, 11, 8, 9, -13, 55, -23, -6, -8, -19, 6, 25, 2, -44, -23, -15, -31, 4, -6, 2, 9, -3, -14, -13, 0, 4, 12, 11, -10, 18, -10, -5, -21, 5, -2, 12, -45, -1, 28, 22, 1, -17, 21, 5, 11, -27, -25, 10, 4, -17, 5, 7, -55, 28, 1, 4, -1, 25, 11, 33, -40, 3, 16, 26, -10, 4, 5, 5, 16, 4, -25, 28, 3, -19, -6, 18, -36, 52, -24, 8, -5, 30, 14, 32, -30, 4, -2, 6, -4, 15, -18, -8, 27, 9, -22, 22, 11, -1, -8, 12, -16, 25, -22, -20, -36, -22, 42, -41, 10, -35, 7, 10, -5, -14, 38, -3, 19, -12, -21, -7, 2, -7, 37, -21, -44, -12, -37, -27, -38, -12, 51, -34, -11, -38, 22, 20, -27, -22, 45, 23, 28, -26, -38, 16, 2, -30, 14, 4, -34, 4, 1, -11, -22, 2, 18, -20, -21, -28, 29, 12, -32, -7, 14, 47, -9, -25, -49, -3, -14, -33, -10, -4, -11, 15, 0, -3),
    (8, 12, -5, 3, 8, -34, 34, 4, 19, -12, -31, -27, -58, 7, -17, 30, 4, 15, -29, 6, -5, 11, 25, 18, -31, 15, -24, -26, 15, 30, -11, -5, -9, -31, 3, 12, -22, -26, -17, -14, -34, -20, -11, -1, 8, -35, 2, 11, 0, 6, -11, -5, -8, 12, -11, -20, -15, -2, 20, -1, -13, 30, 6, -21, 0, 32, 15, 4, -6, -40, -30, 20, 12, 26, 3, 15, 10, -24, 17, 18, 4, -8, -32, 17, -26, 16, -32, 40, 6, 28, -10, 18, 20, -27, 11, 31, -19, 0, -25, 9, 8, 34, -4, 14, 0, -17, 0, -13, 3, -15, -26, -17, -15, -10, 1, 0, -5, -24, 6, -30, 1, -10, 14, -23, -20, 7, -27, 8, 1, 4, 16, -8, -4, 20, 3, -23, 11, 19, 14, -7, 12, 14, -18, 40, 7, 9, -12, 23, 19, -22, 8, -16, -6, -28, -12, 24, -12, 12, -13, 10, 20, 0, 4, 7, 22, -5, 12, 18, -14, 10, -22, 28, 6, -14, 5, 22, 8, 12, 12, -26, -2, 3, -22, 20, -16, 3, -25, 3, -3, -5, 29, -10, -26, 19, -22, -22, -4, 4, -15, -16, -13, 3, 5, -17, 4, 21, -11, 1, -5, -37, -1, -10, -21, 10, 1, -26, -5),
    (-4, 6, -11, -7, 14, 21, 20, 6, 18, 9, 12, -14, -50, -12, -5, 39, 6, 4, 22, -4, -25, 1, 3, 12, 8, 3, 12, -29, -3, 10, 33, -27, -2, 29, 13, -28, -17, 9, 29, -4, -3, -8, -20, 9, -19, 12, 0, -25, -9, 8, -20, -10, -28, -2, 29, -14, 1, -32, -12, 11, -20, -6, -3, -23, 13, -20, -23, 0, -34, -5, -17, 23, 14, 1, 0, 3, 27, 16, -11, -2, 19, 35, 28, -4, -27, -33, -5, -8, -4, -5, 3, -14, -12, 21, -11, -6, 6, 7, -1, 4, -16, 10, 33, 4, 1, -42, -25, 3, 6, -16, -28, 7, 21, 17, -23, 27, -45, 24, -17, -3, -10, 4, -18, -33, 26, -19, -3, -17, 10, -17, 18, 17, 14, -4, -5, -34, 29, -31, -8, -17, 3, -34, -22, 16, 22, 4, -15, 7, -16, 22, -2, 0, -12, 15, -36, 0, -12, -23, -20, -36, -1, 19, -16, -24, 12, 9, -4, -27, -28, 35, -11, 13, -24, 2, -37, 14, 8, -28, -18, -11, 10, -1, -9, 16, 14, -12, -4, 17, -18, 8, 8, 13, 18, -1, -23, -19, 36, 4, -20, -10, -28, 3, 18, 5, -1, -10, -32, -3, 6, 5, -14, -26, 13, -39, 3, -18, -4),
    (-9, 7, -14, -1, -15, -14, 14, -20, -2, 5, 5, -30, -35, 5, -27, 11, 5, -43, -31, -16, -12, 13, 14, 1, -18, 16, 4, -38, -8, -18, 32, -19, 7, -13, -34, 2, -49, -58, -8, 14, -20, -24, -9, -23, -17, 11, -1, -11, -10, 3, 19, -38, -19, -14, 15, -24, -5, 26, 3, -16, -36, 24, -8, 18, 12, 5, -8, 2, 8, 7, -17, -12, 29, 6, 7, -5, -37, -8, 21, -3, 2, -8, 21, -20, -7, 28, 43, -11, 17, -19, -27, 5, 29, 29, 15, -1, 11, 17, -25, -17, 0, -37, 43, -7, 19, -12, 12, -5, -13, 31, 11, -12, 18, -16, -35, 13, 23, 17, 8, 21, 3, 3, -30, -28, -24, -17, 11, -16, -1, -8, 0, 18, 6, -18, -13, 22, -17, 13, -25, -4, -19, -7, 10, 6, 9, -23, 11, -14, -22, 7, 12, 3, -17, -7, 12, 3, 17, 11, 24, -41, 18, -6, 5, -15, -1, -2, -8, 13, 14, -4, -14, 13, -4, -16, 30, -1, 8, -17, 19, 13, -22, 20, 25, -47, 39, 7, -2, 5, 4, -14, 18, 27, 14, -9, -2, 15, 22, -10, 20, -4, 6, -13, -11, 2, -29, 24, -6, 13, 12, 22, -17, -4, 13, -6, 26, 8, 25),
    (-20, -14, -15, -69, -16, 25, -28, 0, 34, -15, -9, 23, -20, -2, -38, 18, -25, -29, -5, 7, -26, -28, 28, -28, 4, -29, -5, -59, 10, 12, -14, 34, 23, -26, 36, -12, 20, 13, 5, -1, -8, 3, -6, -10, -2, 4, -3, -14, 24, -14, 8, -8, -4, -14, 15, 2, -23, -6, 15, -10, 4, 18, 8, -5, 26, 5, -6, -12, 0, 22, 15, 21, -12, -23, -13, -47, -3, 36, 22, 45, 28, -17, 30, 12, 10, -8, -20, 7, -11, -7, 3, -16, -49, -11, 36, -17, 61, -25, -10, -40, 14, 26, 31, 24, -5, 5, 60, -36, 0, -2, 13, 23, 13, 4, -9, -20, -5, 49, 15, -13, 10, -4, -10, 1, 7, -30, 25, -44, -24, 12, 4, 5, -34, -9, 16, 26, 15, -21, -21, 0, 0, 31, -13, 9, 16, 10, 3, -17, 12, 37, -20, 27, -28, -14, 32, -28, 6, -4, -8, 19, -7, 7, 1, 3, 4, 3, 7, -10, 28, -10, 14, -14, 3, 1, -5, 1, -46, -2, 25, -15, -10, -12, -4, 5, 21, -23, -16, -3, 4, 22, 2, -8, -12, -4, -1, -7, -21, -6, 2, -52, -5, -12, -33, 21, -6, -7, 9, -5, 7, -8, -5, 3, 18, -11, -24, 0, -11),
    (13, 8, -11, -10, -13, -12, -9, -15, -7, 11, -3, -18, -31, 13, -8, 21, 20, -13, -17, 37, 9, 4, -5, -3, 3, 13, 7, 46, -21, -29, -11, -22, -8, 15, -20, 27, -28, 10, 9, 17, 11, 2, 16, 19, 4, -8, -30, -5, 12, 3, 19, 40, 2, -10, -1, 3, 0, 21, -18, 14, -9, 3, 12, 4, -17, 6, 29, 4, 7, -11, -16, 18, 36, 4, -7, 2, -16, -21, 29, -12, -10, 18, -10, -8, -57, 27, 6, 11, 48, -14, -20, 38, 0, 29, -4, -16, -4, 14, -10, 29, -38, -21, -6, -23, -23, 29, -34, 22, -30, 13, 31, 14, 28, 1, -2, 45, -4, 4, -52, -12, -4, 26, 12, 31, -19, 5, -27, -5, -5, 20, -30, 20, -3, 12, 19, 6, -1, 12, 20, 28, 1, -13, -33, -3, 33, -6, 2, 1, -28, -5, 27, 5, 3, 2, 3, -12, -31, 22, 11, -6, 37, -5, -23, 22, -12, 8, -9, -5, -12, 6, 8, 10, -30, 4, -14, -2, 7, 21, -13, 19, -20, 7, 12, -19, 26, 2, 8, 22, -13, 3, -27, -3, -4, 4, 16, 19, -21, 10, -34, -3, 12, 6, -13, 11, 13, -2, 20, -5, -9, 3, 29, 5, 4, 2, -11, -22, 3),
    (20, 12, -21, -10, -22, 27, -12, -30, -17, -24, 3, -9, 16, 5, 3, -5, -6, -9, 17, 6, 6, 29, -37, -9, -6, 12, -34, 15, -3, 31, -49, -21, -17, -30, -31, 5, 3, -41, -41, 6, -29, -7, 4, 3, 5, -20, -21, -4, -21, 13, -35, 11, -8, 14, -26, 0, -2, -42, -36, 3, 6, -45, -34, 38, 0, -14, -29, -36, -20, 7, -10, 15, 16, 30, 16, -5, 24, -18, 36, -36, -10, 10, 2, -31, -13, 7, 14, 13, 2, 12, 11, 4, -4, 29, 34, -3, 13, 31, 30, 8, 43, -7, 25, -26, -25, 20, 8, -29, -28, -6, 13, 19, -28, 29, 35, 3, 8, -14, 63, -15, 0, 9, -8, 3, 25, 22, 10, -5, -15, -3, 13, -12, 1, -34, 14, 34, -44, 14, 5, -36, 12, -6, 32, -18, -1, -36, -34, -2, 0, -22, -7, -3, -6, -7, -29, 9, -14, -20, -7, -20, 27, -11, -20, 5, 8, -11, 4, 11, -13, -3, 8, 10, 20, -25, -15, 4, 3, -10, -25, -6, 4, -2, -5, -19, 26, 12, 2, -4, 13, -18, 31, 4, -7, 2, 8, -12, 13, 7, 20, 0, -10, -11, 7, -25, 12, 1, 6, -18, 0, 10, -2, -35, 6, -10, 27, -21, -3),
    (19, -22, 21, -8, 8, 31, -32, 9, -5, 4, 30, -29, 17, -11, 26, -4, -3, 4, 12, -15, -5, 38, -5, -29, 20, -19, 14, -47, -13, 35, -12, -3, 2, -4, 52, -48, 7, -18, 20, -17, 12, -10, -18, -19, -9, 44, 31, -52, 15, -31, -32, -25, -18, -12, 12, -22, 11, -5, 2, -2, 3, 10, 15, -13, 9, -29, -20, 0, 2, 21, 12, -29, 32, -9, 30, -19, 4, 11, -26, 20, -7, 4, 29, -29, -21, -7, 18, -21, -21, 25, -12, -27, -3, 35, -21, -28, 32, -20, 7, -40, -14, -7, -29, -12, -21, -13, 37, -46, -38, -21, 28, -22, -18, -2, -37, -13, 12, 36, 2, -37, 15, 3, -2, -9, -19, -16, 21, 2, -2, -10, -22, -1, -48, 8, -5, -36, 20, 9, -24, 6, -15, 13, 4, 22, 9, 10, 28, 4, 8, 13, -4, 5, -2, 19, 16, -4, -14, 1, 12, -16, 2, 3, -3, -5, 2, 10, -12, 6, 23, -8, 7, 1, -19, -1, -1, -26, 3, -5, 19, 5, -18, 0, 18, -36, 9, 14, -19, 5, -1, 13, -1, -16, 14, 12, -11, 18, -13, -10, 6, 28, 1, -12, 2, 11, -11, -8, -5, -1, 13, 15, 20, 12, -12, 8, 12, -5, -10),
    (-25, -11, -34, 10, -5, -11, -8, -10, -3, -22, -14, -12, -5, -10, -39, -1, -6, -22, -16, 33, 3, -63, 2, 11, -20, -6, -10, 1, -2, -13, -17, -33, 6, -27, -16, 14, -14, -9, -51, -15, -9, -12, 12, 15, 10, -27, -14, 24, -8, 4, 10, 1, 7, -11, 6, -59, -5, -16, -15, 0, -19, 1, -28, 4, 1, -8, -6, 17, -7, 5, 1, -14, -17, 29, 0, 23, -10, 20, -14, 0, 5, -29, 9, 11, 13, 11, -17, -5, -13, -16, 26, 1, -12, -57, -13, -13, -39, 17, -24, 6, -9, 36, -36, -10, -9, -53, -20, 32, 3, -2, -28, 19, -21, -44, -5, -14, -7, -3, -25, -18, -13, -5, -19, -4, -8, 0, -17, -8, -7, -19, -37, 28, 3, -4, -34, 20, -6, -27, -13, -4, -30, 8, -26, -4, 3, 21, 12, 9, 18, 22, -3, 10, 4, 1, 21, -3, 22, -17, 21, 8, -15, -5, 3, -7, 5, 30, 32, -3, 5, 23, 14, -4, 17, 35, -13, -11, -26, -11, 36, -2, 7, -4, 29, 12, -20, -11, 17, -21, -4, 12, 24, -37, 15, 3, 4, -4, -3, 13, -16, -2, -13, -15, 4, -4, 6, 6, 5, 5, -8, 4, 30, -26, -4, -9, 1, -32, 19),
    (-1, -25, 9, 4, 29, -11, -21, 6, 4, -13, -13, -8, 1, -3, -31, 29, -29, 26, 4, -12, 16, -18, 7, 2, 3, -12, -7, -22, 5, -15, -28, 19, 17, -20, -3, -10, 11, -20, -12, -32, -1, 25, 4, -6, 9, 21, -1, 2, 22, -5, -3, -36, -27, -31, 3, 38, -24, -7, -39, -26, 5, 11, -2, 18, 20, 10, -21, 19, -13, 6, -9, 21, -3, 2, 10, 11, 36, -15, -19, -1, -18, 7, -6, -20, -13, 11, -21, 16, -30, 36, 8, -1, 22, -26, 2, 3, 25, -12, 14, -4, 43, 1, -3, 17, -7, -11, 33, -21, -25, -22, -24, -61, -19, 18, -2, -39, -1, -3, 1, 3, 18, -5, 13, -27, -15, 12, -19, 35, -24, -20, -39, -24, -12, 9, -12, 41, 29, -3, -32, 26, 12, 12, 6, 16, -7, -4, 7, 14, 20, -20, -14, -1, 8, 24, -12, -1, -13, -16, -5, -4, -7, -1, -1, -10, 10, -12, -11, -16, 12, -17, 1, 8, 6, -45, -23, -13, -27, -15, -21, 4, -6, -36, -16, -58, -38, 20, -25, -33, -1, -9, -17, -15, 44, -20, -4, -10, -14, 13, 5, 20, -18, -24, -27, -18, 11, 32, -15, 32, 3, 4, 4, 27, -18, 18, 1, 9, -5),
    (25, -17, -13, 14, -25, 12, -22, -3, -21, -3, 5, -9, 17, 6, 12, -16, -9, 5, 15, -14, 22, 20, -25, -2, 35, -15, -18, 28, -6, -41, -22, -4, 2, 18, 6, -2, -7, -16, 3, -31, -9, 32, 0, -7, 20, -6, -26, 17, 20, 19, -9, 33, 26, 9, 16, 6, 3, -22, -31, 35, -32, -12, -43, -13, -10, 14, 6, 10, -12, 9, -19, 18, 17, -5, -10, 1, -15, 11, -17, -19, -56, 11, 11, -18, 7, -13, 22, 20, -10, 13, 13, 10, 3, 38, -11, -27, -4, 1, 1, 20, -5, -19, -4, -65, -39, 49, -27, 21, -31, -8, 21, -23, -11, -2, 8, 27, 11, 24, -36, 9, -20, 29, -16, 31, -12, 51, -32, 0, 17, -21, -7, 24, 12, -19, -26, -19, -48, 22, 36, -19, -28, -33, -62, 6, 9, -6, 16, 13, 12, -4, 4, -11, -36, 26, 0, 19, -4, -8, 18, 2, 12, -11, -2, 18, 7, 4, 25, -11, -18, -4, 12, 26, -41, -16, 7, -44, 4, -15, -41, 33, -12, -50, -3, -40, -6, -26, 15, -9, -24, -14, -15, -8, -25, 2, -23, 30, 4, 36, -12, 34, 24, -29, 17, -22, 27, -3, -34, 3, -4, 1, 12, 15, -30, -17, 24, -27, -22),
    (-4, -31, 23, 3, 13, -30, 5, -1, -1, -5, -13, -3, -15, 2, 0, -9, -5, 12, 8, -4, 27, -13, 16, 0, 5, -30, 28, -13, 23, -28, 3, -3, -15, -21, -3, -13, -20, 5, -13, 17, 9, 11, -9, 11, 42, -36, 4, -3, 2, -10, 18, -8, 0, -38, -2, 1, -6, 4, -13, 5, 1, -5, -11, -22, 8, 3, -13, -4, 20, -13, 17, 1, 3, -48, 20, 23, 17, -24, -32, -12, -24, 8, -22, 7, -4, 4, -4, 9, -6, 10, 4, -12, 30, -31, -29, -28, 11, -57, 13, 14, 32, -67, -52, 2, -7, -4, -21, -13, -12, 8, -24, 15, 1, 8, 4, -3, 36, -45, -28, -6, 3, 4, 2, 7, 5, -30, -8, -7, 16, 7, -2, -3, 20, -50, -35, -39, -16, 7, -6, -29, 29, -21, -15, -5, -6, 1, 21, 3, 2, 6, -29, -13, -17, 8, -6, 17, 2, -2, -4, 11, 2, -3, 3, -4, 20, -20, -21, -13, -13, 0, 20, -2, 7, -36, -43, 0, 12, 11, -5, 5, -7, 0, -7, -25, -19, -6, 14, -4, 33, -15, -35, -24, 4, 3, 0, 9, 8, -29, -3, -25, -4, -12, -20, -12, -5, -39, 4, -35, -43, -10, -3, -16, 20, -9, -27, 2, -9),
    (5, -1, 4, -16, -4, -25, -2, 12, 15, 4, -12, -26, -33, 4, -14, 21, 22, 12, -33, 6, -21, 11, 3, -24, 17, 1, -2, -9, -5, -22, 14, -21, -24, 30, -15, -8, -19, 13, 4, 42, 20, -11, -14, 34, 18, 29, -6, -11, 12, 26, -1, 11, -12, -19, 19, -29, -35, 20, -20, -6, -17, 22, 15, -6, 23, -2, 12, 9, -5, 0, -21, 6, -11, -7, 4, 19, -3, -10, 12, -8, 29, 5, 1, 15, -8, -3, -22, 21, 0, 22, -14, 28, -27, -22, 22, -21, 31, -16, -20, 30, -17, -39, 24, -13, -2, 23, -23, 4, -48, 28, 0, 17, 44, 10, -16, 31, 3, 20, -4, -1, 3, -8, 3, 2, -18, -38, 11, -12, -36, 21, -37, 1, -33, 7, 29, -13, 11, 12, 13, 21, 3, 7, -35, 29, 3, 17, -9, 38, 6, -32, 19, 11, 19, 5, -4, 19, -2, -2, -2, 24, 15, -6, -12, 8, -39, -13, 1, -7, 17, -1, -23, 19, -26, -28, 24, -11, -13, -4, -11, -13, -48, 11, 10, 6, 23, 3, -17, 23, -7, 6, -16, 27, -13, -8, 12, -13, -1, -1, -6, -6, -36, 12, -25, 11, 0, 10, 10, 4, 4, 12, 19, -4, 5, -12, -23, 31, 23),
    (7, -12, -1, 22, -9, -38, 1, 6, 13, -7, -28, 21, -6, -20, -25, -28, -17, 29, -16, -1, -11, -12, -6, 17, -10, -6, -21, 19, 18, 1, -12, -12, 9, -37, -18, -10, -13, 8, -38, 10, -14, -11, 4, 8, -33, -8, -25, 3, -37, 16, -19, 14, 11, 10, -19, -11, 16, -33, 6, 1, -9, -20, -46, -17, -17, -38, 12, -3, -17, -25, -9, 25, -47, -21, -27, 4, -27, 2, 18, -18, 3, -15, -4, 5, -15, 10, 2, -27, 7, -21, -12, 2, -7, -39, 0, -6, 8, -5, -13, -20, -18, 1, 6, 35, 3, -23, 2, 10, 5, 4, -4, -9, -30, 1, 11, -8, -34, 7, 10, 2, -24, -17, -29, -13, -13, -17, -6, 33, -6, -15, 11, -29, 28, -11, 4, -6, -29, -6, 4, -38, 3, -31, 0, -3, -8, -6, -11, -12, -13, 44, 11, 29, -7, -33, 12, 8, 49, 12, 19, -29, 14, -26, 20, -5, 11, -5, 27, -22, -19, 4, -8, -28, -2, 36, 0, 38, 12, -11, 19, -16, 39, -9, 6, 16, 12, -31, 4, -6, -6, 43, 13, -48, -4, -12, -1, -21, 1, -9, 29, -6, -18, 10, 4, -11, 11, 3, 17, -2, -15, -20, -3, -29, 7, 36, 5, 1, 33),
    (-21, 1, -4, -4, -12, 17, -11, -1, -27, 3, 4, -13, 10, -8, -12, 3, -16, 19, 23, 29, 12, -14, -18, -8, -6, -12, -9, 6, -12, 20, -48, -4, -42, 4, 4, -21, 12, 2, -4, -21, -20, 4, 26, 22, 14, 4, -32, -19, 10, -7, -29, 11, -1, 1, -30, -24, -21, -3, -11, -4, 4, -9, 3, -34, -24, 4, 4, -2, 9, -29, -13, -6, 3, -3, 19, -16, 0, 33, 28, 19, 0, -4, 27, -41, 21, -30, 12, -1, -29, 29, 23, -22, -23, 30, 20, -29, 31, -9, 12, -49, 5, 55, 43, 22, -36, 10, 56, -73, 12, 9, 38, -28, -23, 12, 23, -34, -36, 66, 11, -43, 30, -6, -12, -34, 19, 42, 17, -1, -24, 9, 21, -20, 3, 22, 20, -31, -16, -4, 7, 2, -4, 33, 14, -20, 5, 12, 4, -26, 10, -4, 5, 18, 8, -15, 5, -21, 11, -11, -13, -5, 2, -5, -23, 3, -6, -10, 11, 8, 24, -15, 16, -14, -10, -26, 14, 11, 1, 2, 19, 1, -12, 23, 0, -7, 7, 1, -45, 12, -9, 24, 2, 27, 12, -27, -4, -8, -23, 3, 17, -31, -5, 10, 11, 13, -11, 21, 1, -9, 19, 13, -38, 2, -12, 20, 22, 30, -7),
    (13, -25, -14, 0, -19, 8, -12, -17, -3, -5, 19, -1, -46, 26, -8, -25, 1, -32, -7, 16, -13, -21, -21, -17, -4, -2, 17, 29, -4, -2, -27, -4, 9, -10, -10, 23, 20, 41, -14, -11, 23, -10, 14, 14, -6, -6, -58, -2, 4, -18, 22, 5, 3, 14, 3, -17, 25, -12, -4, -2, 28, 23, 0, -10, 23, -2, -5, 21, -11, 8, -7, -1, 12, -8, -5, -33, -36, 15, 26, 3, -15, 12, 14, -2, -12, 21, 2, 6, 13, 8, 7, 1, -35, -5, -9, -10, 24, 14, -14, 35, -23, 22, -20, 5, 19, 6, 13, 17, 12, 49, 20, 10, 9, -1, 10, -5, -89, 20, -60, -4, 11, 14, -12, 14, -21, 20, -21, 4, 28, -8, 1, 21, 20, 20, 13, -29, 1, -15, 15, 4, -63, 32, -49, 13, 19, -1, -9, 5, -29, 22, 10, 3, -33, 7, 13, 6, -10, 6, 16, 8, -3, 6, 3, -1, -47, 16, -11, -10, 33, -6, -17, 18, -39, 19, -19, 4, -11, -3, 7, 0, -2, 7, 16, 4, -10, 1, 6, -6, -50, 23, -21, -10, 14, 2, -19, -11, -36, 10, 1, -1, 11, -1, 8, -9, 3, -37, 5, -19, 11, -12, 3, -23, -28, 13, -8, -10, 49),
    (-46, -14, -14, -31, -13, -15, 6, -51, -21, -15, -25, 10, 7, -12, -22, -21, 3, -56, 3, 26, 4, -26, 2, -7, -17, 2, -21, -15, -13, -23, 5, -8, -24, -37, -33, -32, -16, -13, -4, 27, 5, -7, -29, 13, -2, -22, 25, 29, -9, 17, -5, -18, 27, -8, -16, -4, 3, -12, -11, 9, -24, -3, -19, 22, 2, 3, -10, 8, -5, -29, 5, 16, -9, 4, -11, -30, -2, -19, 42, 29, 22, -15, -8, 14, -57, 23, -12, 3, 20, 4, -34, 15, -6, 7, 50, 14, 10, 12, 10, 14, 16, -12, 23, 13, -20, 10, -22, 11, -25, 4, -29, 52, 18, 13, -36, 5, -4, -2, 24, 20, 20, 12, -10, 10, 32, 3, 1, -9, -19, 14, -14, 13, -27, -29, -29, 52, 8, -3, -29, 12, -11, 14, 6, -9, 6, 6, -12, 27, 8, -4, 11, 24, 16, -11, 4, 14, -11, 6, -18, -6, 12, 11, -4, 23, 9, -9, 16, 37, 23, 5, 2, 9, 8, -37, 13, 31, 20, 1, -9, 5, -15, 5, -39, 30, 16, 24, -41, 33, 11, -7, 26, 44, 11, 11, -10, 6, 22, -12, 10, -9, -2, 16, -11, 4, -20, -29, 0, 8, 16, 4, -36, 19, -7, 10, 20, 23, 37),
    (2, -40, -4, -10, 13, -4, 15, 22, 11, 10, 3, 1, 29, 4, -27, -16, -10, -24, 15, -20, -14, 5, 36, -48, 20, -30, 19, -38, 6, -17, 30, 5, -28, 18, 2, -30, -7, 5, 19, -35, 20, -9, -6, -34, 12, 4, 19, -11, 12, -21, 12, -12, 4, -17, 35, 5, -11, 0, 10, -13, -20, 2, 11, -33, 18, 3, -15, 14, 22, 2, 18, -1, 21, -4, 15, -50, 12, -4, 4, 18, -5, 3, 14, -7, -13, 22, 18, 31, 30, 2, -14, 21, -13, -39, -6, 1, -5, -35, 15, 8, -14, -12, 13, -5, 17, 24, 9, 8, 7, 23, 12, -29, 38, -6, -6, 18, 1, -16, -19, -21, -5, -13, 18, 14, -10, -5, 5, 4, 34, 4, -4, 3, 6, 10, 12, -60, -4, 12, -1, 14, 22, -5, 5, -28, 18, -11, -5, 14, 5, -12, -37, -18, -19, 2, -5, -19, 4, -29, -3, 12, -20, 16, 15, 18, -4, 19, -11, 8, 12, -17, 26, 20, 6, 13, -37, -3, 2, 20, -2, 2, 3, -7, -25, -3, 1, 4, 17, 8, -4, 0, 3, 4, -25, 3, 19, 1, -1, 5, 1, 11, 12, -4, 6, -13, 2, 25, -2, -14, 23, -9, 20, 14, 11, -14, 5, -13, -16),
    (5, -6, 13, -24, 16, -13, 29, -13, -18, 23, 13, -9, 1, 15, 23, 13, -2, -62, 5, 13, -26, 28, 10, 16, 6, 13, -21, -9, -10, -1, -5, -81, -10, -4, 4, 1, 23, 0, 27, 29, 0, -60, 14, 20, -14, 11, -26, 20, -5, -15, -17, 22, -20, 18, -22, 0, 11, -7, -9, 3, 36, 29, 3, -11, -3, 6, 1, -3, 4, 14, -6, 4, -23, 31, -10, -22, -18, 23, 21, 12, -16, -9, -4, 15, -26, -18, -58, 4, 5, -3, 1, -4, -37, -20, 28, 13, -18, 14, 0, -18, -33, 20, -16, -15, 20, -7, -3, -2, 9, -29, -18, 1, -23, 1, -3, -29, -51, -12, 9, 2, -5, -39, -21, 31, -37, -17, 2, 19, -6, 5, 3, 3, -32, 38, -13, 6, 30, 0, -8, 28, 9, -19, -21, 20, -5, 27, -16, -2, 25, 17, -12, 2, -14, 5, 12, -8, -1, -13, -11, -1, -35, 9, 26, 6, 1, -16, 12, -12, -8, 36, -6, -3, 23, -4, 13, 6, 1, 9, 19, -6, -9, -28, -16, 12, -29, 6, 11, -15, -12, 6, 10, -5, 9, -27, 3, 8, -15, -31, 10, 9, -12, 0, 7, -3, -29, 22, -8, -6, 27, 8, 2, 30, -22, 10, 2, 14, 0),
    (13, 4, -23, 0, 5, -15, 11, -59, 20, -46, -39, -27, -26, -11, -10, -55, 11, -7, -13, 0, -26, 26, -52, 19, -14, -13, -20, 11, 5, 5, -21, -11, -2, -35, -32, 4, -17, -6, -65, 33, -19, 1, -15, 30, 0, -16, -11, 10, -43, -19, -16, 10, 27, -25, -34, -3, -4, -12, -27, -3, 10, -2, -40, 6, -28, -7, 5, 10, 30, -45, 4, -5, 5, 16, 14, -4, -3, -23, 2, -17, 5, -28, -28, 18, -29, -14, 5, -23, -13, -25, -13, -15, -29, 20, 3, -6, -16, -5, -12, -4, 15, 36, -26, 20, 4, -17, -7, 29, 19, 3, -49, -6, -32, 2, 2, -4, -21, -12, -4, -6, 24, -11, 12, -9, 20, -5, 3, 23, 1, -10, 7, 8, 21, 20, -15, 6, -5, 14, 17, -12, -8, 24, 4, 20, 25, -1, 11, -10, -18, -23, -17, -21, -3, -14, -17, 14, -26, 8, -1, -20, 7, -9, -20, -7, -29, 16, 5, -13, 20, -3, 0, 7, 2, 36, -1, 16, 2, -30, 22, 9, 28, 0, -15, -11, -15, -19, 9, -4, -41, 31, -4, -4, 37, 1, 24, 3, 17, 5, 22, 15, 6, 3, 13, -1, 5, 11, 4, 14, 6, 15, 11, -19, -20, 11, -12, 3, -2),
    (-15, 17, -13, 18, -42, 15, -2, 26, -20, 4, 15, 23, 23, 23, 18, 14, -18, 11, 4, -13, -32, -6, -6, -2, 7, 4, 21, 13, -36, 12, -15, 40, 7, 6, -1, 15, 13, 18, 2, 18, 7, 17, 8, -27, -67, -13, -23, 11, 5, 19, 9, -3, -8, 20, -1, 40, 14, 5, -16, 6, 13, 13, -6, 7, -4, 1, 2, -29, -34, 1, -1, 27, -9, -9, -19, -8, -50, -3, -21, 3, -27, -13, 14, -6, 13, -18, 23, 4, -3, 9, 3, 1, -16, 17, 7, -27, -2, -17, -6, 0, -30, -14, -18, 17, 3, -9, -15, 0, -10, 0, -7, 19, 10, 12, -1, 1, -33, 8, -7, -18, 6, 8, -17, 2, 9, 27, -17, 20, 9, 4, -4, 9, -9, 10, -12, 20, -31, 11, -1, -3, -54, 16, -2, 17, -2, -2, 2, 22, -4, -30, -1, -45, -20, -25, -15, -7, -2, -29, -3, -1, -21, 20, -7, -32, 33, -4, -1, 14, 12, -41, -4, -19, -12, -45, 1, -5, -3, -40, -7, -11, -3, -19, -15, 6, 20, 12, -19, 8, 15, -20, 29, 18, 3, -14, 6, -15, 12, 16, -4, -6, -5, -7, 2, 15, 7, -14, -30, -5, -10, 15, 12, -6, -21, -11, 3, 10, 45),
    (12, 6, -21, -52, -26, 4, 29, -3, 14, -25, 20, -24, -23, 12, 26, 14, 16, -23, -22, 5, -4, -16, 31, 6, 6, 8, -9, -63, -10, 10, 40, -5, -2, 10, 22, -31, -3, 28, 28, 29, 29, -7, -4, 7, 3, 22, 42, 7, 13, -2, -42, -4, -13, 3, 11, -55, -11, 4, 20, -22, -2, 13, 1, -3, -5, -9, -4, 11, -13, 12, 4, -7, 25, -17, 11, 17, -3, 20, 44, 28, 34, -21, 20, -14, -5, 13, 7, -34, 27, 21, -9, -2, 9, -16, -4, 27, 12, -9, 28, 13, -3, -29, 59, 14, 16, -45, 11, -12, -36, 33, 13, -28, 69, 10, -16, -11, 8, -21, 14, 28, -18, 15, 1, -3, 7, -16, 26, -14, -19, -26, -36, -10, -39, 19, 0, 21, 30, -2, -5, -4, 19, -19, -2, 15, 6, -28, -3, 21, -3, 7, -24, 21, 8, 2, -9, 13, 14, -35, -13, -3, -22, 4, 12, -9, -11, -24, 11, -16, -6, -25, -2, 22, -13, -10, -38, 3, -5, -23, -3, 29, 18, -5, -13, 13, -3, 0, 4, -2, 12, -22, -7, 9, -1, -4, -22, 20, -18, -5, -43, 20, -11, -14, -3, 21, 8, -43, -24, 33, -50, 6, 3, -7, -14, -33, 11, -13, -3),
    (20, -17, 3, 3, 5, 5, 3, -2, -45, 21, 16, -35, -11, 13, 17, -4, -17, 28, 7, 3, -3, 12, 12, 33, -4, 0, -9, 4, 7, -31, 35, -35, -44, 22, -15, -13, -19, -30, 7, -27, -13, 24, 0, 4, 8, 13, -12, 50, -12, 6, -25, 10, -16, -7, 6, -13, -1, -8, -11, 11, 12, 27, 3, -7, -4, 8, 17, 12, 1, -27, -6, -15, 4, 2, -19, 3, 13, 2, 38, -13, -38, 18, 10, -17, -13, 11, 11, -56, 13, 21, 15, -14, 5, 11, 5, 52, -4, 26, -25, 20, 21, 3, 20, -48, -28, -36, -28, 5, -12, -30, -19, 13, -45, 29, 4, -3, 13, -9, 17, 63, -9, -10, -19, 30, 3, -17, -22, 13, 5, -30, -16, 29, 18, -19, -22, 13, 20, -3, -6, -5, 20, -61, 18, -46, -4, 20, -12, -4, 3, -13, 19, -28, -2, 9, -4, -28, -4, 9, 4, 0, 8, -3, 1, 9, -4, 13, -10, 34, -6, 16, -13, -9, 10, 11, -16, -42, -2, -42, -4, 35, 11, -19, -19, 54, -30, 19, 14, 3, 16, -12, 4, 5, -16, -14, -14, 4, -1, 9, 2, 3, 28, -3, -8, -3, 26, -13, -5, -7, -9, 9, -15, -10, -27, -13, -5, -36, -15),
    (12, -14, -7, 3, 6, 10, -9, -7, -1, -5, -6, 1, -6, -20, -10, 4, -1, 28, -9, 20, -4, -10, 3, 16, 18, -14, 14, 22, 24, 13, -27, -21, 4, 21, -5, 11, -12, 10, -23, 34, 5, 12, 18, 9, -10, 8, -11, 5, -12, -25, 11, 10, 0, -11, -1, -9, 22, -8, -1, 1, 5, -20, -17, -44, 14, 5, 11, 25, -1, -11, -31, 0, 22, -21, -35, 1, -20, -20, -5, -25, -37, 7, -3, -13, -17, -36, -4, 12, -37, 25, -9, 18, 13, 25, 12, -5, 24, -22, 4, 32, 31, -24, 6, -60, -10, 29, 11, -2, -21, -19, -22, 43, -18, -3, 2, 12, 26, 20, -26, -7, -12, -18, -17, 5, -5, -19, -27, -17, 8, -38, -44, 39, -2, -27, -41, -63, -57, 12, -14, 19, 0, -11, -54, 12, 18, -12, -19, 8, -7, 5, 6, -20, 4, 1, 1, 4, 10, 12, 11, 1, 1, 1, 0, 12, 5, 26, 17, 11, 16, -12, -12, 13, 10, -39, 28, -27, 18, 28, -6, 3, 4, -5, -2, -24, 8, -3, -13, 22, 16, 15, 9, 8, -31, 6, -33, 17, -29, -12, 15, -10, 4, -44, -36, 27, 23, -58, -14, -14, -16, 7, 1, 9, -10, -6, -4, 23, -12),
    (-18, 0, -14, 17, -14, -39, -23, -20, 35, -5, -49, -18, 19, -5, -38, 31, 8, -2, -12, 30, 16, -21, 16, 5, -60, 2, -12, -8, 36, 22, -12, 1, -5, -14, -20, 19, -2, -25, -72, 36, -22, 8, -5, 5, 16, -16, 15, 11, 10, 0, -3, -18, 19, 15, -27, 3, -15, -4, 7, -17, 15, -4, -7, 13, -6, -2, 1, -10, -13, 21, 12, -18, 2, -15, -17, 2, -20, -45, -19, -6, 0, -40, -10, 29, 27, 8, -27, -11, 1, -1, -8, 9, -14, -54, 34, 1, 6, -8, 17, 0, 30, -14, -12, 32, 7, -12, 9, 0, 10, -21, -21, 48, -31, 22, 4, -9, -4, 7, 18, 5, 26, -8, 14, 11, 25, 0, 17, 6, -22, 36, 14, -27, 4, -38, -6, 49, -29, 7, 9, -12, -18, 3, -7, 4, 15, -28, 10, -29, -27, -33, -3, -21, -8, -31, -20, -11, -13, -12, -4, 5, 4, 8, -4, -10, -6, -28, 0, -8, 26, 3, 20, -5, 7, -7, 8, 11, 9, 26, 2, 5, -13, -8, 1, 12, -23, 26, -1, 12, -12, 0, 1, 4, 11, -6, -16, 30, 28, -16, -8, -12, -1, 17, 3, -11, 7, -22, 1, 20, -27, 5, 1, 13, 5, -1, 2, -18, 8),
    (-16, 4, 6, 15, 14, 20, 5, -4, 14, 4, 17, 0, 14, 30, -7, 28, 21, -19, 19, 21, -18, 16, -34, 7, -27, -13, 18, -11, 2, 25, 12, 5, 62, -38, 14, -13, 44, -9, -22, -12, 12, -20, -16, 13, -11, -13, -33, -21, 4, -4, -23, -16, -21, 7, -7, 10, -10, -48, 1, -13, 4, 27, 5, -27, -23, -21, -12, -33, 11, 29, -1, 3, 9, -16, 4, 18, 26, -7, -15, -7, 12, -3, 23, -13, 15, -32, -24, 22, 5, 15, 11, -14, -10, 21, -43, -1, -18, -2, -14, -11, 16, -6, -3, -5, 20, -32, 17, 5, 27, -23, -20, -28, -37, -20, -37, -8, -10, 9, -25, -32, -20, 1, -21, -12, -36, 22, 7, 8, 14, -24, -11, -15, -4, 16, -14, 11, -12, -48, -7, 13, -10, 9, -13, -23, 10, 20, 11, -25, 18, -23, 9, -8, -14, 8, -1, -34, -1, -10, 10, -38, -34, 3, -17, -15, 16, 5, 5, 5, 23, -2, -37, -14, 10, -33, 2, 5, -26, 22, -40, 5, -38, -5, 7, 21, -1, 7, -8, 50, 8, 12, -20, 7, -3, -4, 18, 0, -13, 25, 5, 14, 6, 8, 4, 0, -29, 27, -8, 8, 7, 12, 12, 6, 10, -29, -10, 28, 14),
    (-6, 3, 4, 25, 4, 4, 14, 18, -22, 1, -3, 9, 20, 16, 15, -10, 28, -11, 12, -21, 11, -29, 12, 11, 1, -4, 17, 14, 1, 9, 22, 35, 12, -4, 0, 9, 36, 44, 19, -30, 25, -3, 12, 3, 9, -19, 20, 10, -6, 2, 20, 20, -4, 13, -3, 13, 20, -3, 5, -2, 7, 29, 13, -12, 12, 6, 15, -4, 8, 3, 7, -5, -25, -12, -19, 20, -5, 1, -15, 22, -17, -8, -10, 20, 29, -14, -10, -21, -6, 3, 21, -15, 1, -27, -3, -26, -19, -20, -13, 10, -12, -4, -36, 44, 4, -39, 1, 12, 50, -18, -13, -16, -4, -20, 14, -37, 5, -18, 4, -48, -7, -27, -8, 0, 4, 2, -33, 31, -2, -30, 6, 8, 20, -58, -11, 16, -29, 12, -2, -39, -4, 12, 3, -33, -5, -30, -24, 18, -3, -6, -24, 5, -9, -13, 20, 2, 19, -38, -3, 6, -36, -13, -4, -13, -28, -14, -11, -49, 4, -39, -6, 4, 9, 0, -11, 22, 6, -6, 14, 15, 11, -44, -16, 30, -53, -25, -7, -17, -33, -5, 9, -86, 31, -21, -36, -6, 2, 3, -4, 10, -4, 2, 9, -12, -29, -67, -12, 43, -5, -20, -14, -10, -20, 12, 1, -45, 12),
    (-23, -14, -25, 5, 12, -2, 5, 18, 14, 10, -6, 28, -2, -36, -24, 30, 1, -11, -12, 7, -27, -13, -34, 12, -27, -27, -13, -20, 6, -5, -3, 9, -16, 15, -12, -3, 11, -60, -8, 12, 6, -37, 5, -12, 14, -6, -21, -22, -14, -2, -9, -36, -18, -7, 4, -12, 3, 19, 1, -15, 15, -19, 22, -1, 18, -28, 0, -20, -9, -13, 16, 1, -41, -11, -1, -4, 20, 7, -16, 17, -9, 4, -9, 10, 11, -33, -60, 33, -26, -2, 20, 12, 12, -41, -12, 4, -16, -29, -4, -26, 31, 2, -39, 25, -24, -8, 4, -24, 26, -52, -27, 45, -20, -11, 11, -13, 16, -21, -33, -46, -20, -20, -14, -16, -3, -1, -4, -47, -3, -25, 3, -9, 12, -35, 2, -19, -4, -26, -29, -1, 29, -8, -18, -12, 10, 6, 21, 1, 2, 26, -8, 21, 0, 12, 2, 25, 18, 5, 4, 17, -13, -7, 14, -1, -21, 14, -20, -7, 13, -9, 28, 17, 26, 20, -10, 29, -4, 30, 16, -10, 14, -13, 2, 30, -29, 10, 26, -16, -12, 4, -29, -28, 2, -6, 0, 11, -11, 5, 2, -4, 3, -5, 20, -24, 11, -20, 6, -11, -20, -3, -4, -22, 19, 4, -23, -38, -2),
    (-33, -1, -24, -46, -4, 27, -21, -28, 0, -27, 3, -6, -35, 2, -19, 5, 4, -20, -20, 11, -20, -22, -46, -11, -60, 6, -12, -6, -4, 4, -23, -13, -11, -39, 3, 18, -8, -4, -8, -26, -19, -40, 13, -31, -24, -16, -34, -11, -22, 10, -20, -10, 0, -22, -11, -7, -6, -27, -4, 10, -21, 5, -10, -16, -13, -29, -2, -22, -39, 8, -8, 0, -12, 16, 15, -22, 27, 17, -8, 16, -29, -13, 13, -12, 23, -24, 28, 29, -5, -34, 6, -22, -1, 11, 31, -21, -1, 23, -4, -33, -4, 31, -17, 17, -24, -16, 16, -27, 23, -44, 31, 20, -20, -34, 5, -30, -12, 33, -4, -23, 12, 23, -5, -12, -19, 16, -14, 12, -31, -24, -7, 9, 6, -16, 13, -24, -5, -3, 4, -15, 11, 17, -25, -12, 5, 26, 20, 11, 20, -3, 5, 17, -9, -6, -10, 5, 12, -37, -13, 36, -20, 4, -4, -4, -7, 1, 16, 10, 3, 40, 27, -22, 10, -4, 28, 10, -17, 6, -5, -8, 22, -41, -3, 29, -20, -15, -5, -9, 21, 5, 26, 14, 4, 11, 11, -11, -4, -5, 5, -12, -7, 23, 12, -6, 4, -2, 6, -6, -7, -12, 2, 1, 27, 4, 5, 14, 2)
  );
  ----------------
  CONSTANT Layer_6_Columns    : NATURAL := 4;
  CONSTANT Layer_6_Rows       : NATURAL := 4;
  CONSTANT Layer_6_Strides    : NATURAL := 2;
  CONSTANT Layer_6_Activation : Activation_T := relu;
  CONSTANT Layer_6_Padding    : Padding_T := same;
  CONSTANT Layer_6_Values     : NATURAL := 32;
  CONSTANT Layer_6_Filter_X   : NATURAL := 3;
  CONSTANT Layer_6_Filter_Y   : NATURAL := 3;
  CONSTANT Layer_6_Filters    : NATURAL := 32;
  CONSTANT Layer_6_Inputs     : NATURAL := 289;
  CONSTANT Layer_6_Out_Offset : INTEGER := 6;
  CONSTANT Layer_6_Offset     : INTEGER := 0;
  CONSTANT Layer_6 : CNN_Weights_T(0 to Layer_6_Filters-1, 0 to Layer_6_Inputs-1) :=
  (
    (21, -15, 22, 10, -12, 35, -9, 4, -8, 5, -4, 0, 36, 19, 20, -10, -14, 3, -4, -8, -9, -2, 33, 1, -26, -17, 12, -3, 22, -27, -17, -18, 7, -12, 28, -8, -17, 23, -2, -7, -20, -22, 3, -19, 35, -21, 22, -17, -11, -1, 0, -3, 5, -3, 19, -15, -6, -8, 2, 32, 28, -20, 23, -20, -3, -16, 28, -18, -12, -3, 1, 3, -14, -26, 10, 13, 10, -2, 8, 4, -1, 12, -23, -2, 23, -28, 9, 0, -6, -8, 1, 15, 24, -11, 19, -15, 14, -35, -3, 30, -13, -5, -6, 1, 7, -8, -3, -8, -6, -9, 19, -18, -4, 11, -1, -23, 0, 32, 15, 4, -31, 9, 30, -24, 11, -24, -13, -25, 21, -4, 45, -8, -17, 20, -38, 7, -6, 2, 12, -45, 25, 3, 3, -38, -29, 12, -21, -6, -4, -14, 19, -10, -14, -9, 20, -6, 4, -30, 11, -30, 15, 4, -4, -22, 6, 15, -8, -48, -12, -11, 0, 11, -14, -11, 7, -8, 12, -13, -16, -14, -15, -12, 3, -26, -17, 10, 5, -6, 18, -2, 14, -2, -21, -4, -8, -10, 21, 2, -11, 4, 19, -24, -11, -19, -21, 44, 2, -2, -9, 4, -2, -10, 12, 11, -5, -11, 13, 28, -3, -12, -9, -3, -17, -13, 22, 3, 13, 24, 1, -5, -7, -22, 5, 20, 5, -5, 12, -11, 18, -24, 16, -2, 7, 18, 2, -7, 7, -5, -19, 3, 18, -17, 0, -20, -16, -21, 16, 13, 3, 1, 16, 0, 26, -20, -12, 1, 21, -5, 24, -19, -6, -14, 1, 7, 25, 20, -14, -7, -6, 18, -6, 29, 3, -10, -5, -27, 2, 16, -8),
    (7, -1, 12, 11, -4, -2, -24, 1, -7, 3, -17, 14, 26, 0, -24, -14, 12, 9, -8, -12, -11, 3, 30, 12, -12, -3, -11, -2, 30, 1, 15, 19, 2, 2, 22, -35, -14, -5, -5, 3, -7, -23, 4, 12, 16, 7, -30, -4, 20, 28, -6, -2, -10, 0, 24, 15, 3, -5, -31, 5, -11, -1, 9, -10, -5, 4, 28, -20, 7, 12, 25, 19, -10, -11, 26, -7, -8, 4, -18, 17, 9, 2, 6, 4, 0, -1, 13, 0, 8, 12, -12, -30, -5, -5, 16, -6, 3, 0, 13, -4, -17, -7, -27, 29, 4, -20, -3, 37, 21, 15, -4, -4, 8, 20, -4, -1, -12, -13, 29, 1, 9, -20, 24, 21, 28, 10, -15, 6, -7, 0, 21, -25, -12, 12, -20, 20, 12, -18, 5, 20, -14, 5, -36, -8, -1, 13, 2, -1, -5, -9, 46, 3, -6, -7, 29, 25, 28, 0, 6, 2, 2, -2, 15, -9, -21, -3, 9, 23, -6, -20, -4, 17, -27, 6, -40, -5, 17, 10, 1, 3, -11, 3, -9, -20, 18, -8, -29, 18, 16, -7, 19, 18, 2, -22, 2, 2, -19, -11, 11, 23, -4, -14, 12, -10, 3, 26, 9, 18, 12, -1, 8, 2, -4, 6, 13, -12, 20, -17, 3, -4, 9, 13, 4, 24, -4, -12, 13, -13, 22, 4, 24, 19, 5, -47, 7, -5, -23, 1, -17, 5, 6, 5, 8, 5, -19, -6, 17, 12, 26, 15, 27, 13, 37, -3, 12, 14, -3, -3, 11, -11, 3, 7, 16, 0, -20, -31, -3, 6, -9, 0, -35, -28, 34, -7, 14, 22, -33, 7, 6, 1, 30, -29, 13, 3, 13, -4, 15, 10, 19),
    (-12, -20, 6, -13, -9, -15, -19, -3, -6, -36, 9, -11, -14, 14, -26, -8, -7, 13, -1, 14, -16, -22, 19, 5, 20, -15, -19, -26, 16, 5, -3, -6, -24, 7, 4, 16, -2, 0, 2, 12, -20, -19, -10, 14, 18, 26, -14, -13, -12, -5, 18, 6, -34, -1, 30, -11, 24, 4, 21, -5, -6, -4, 8, -15, -13, 10, -10, 11, 10, 19, -3, 26, -19, -21, 9, 13, 25, 0, -14, -22, 6, -21, -2, 13, -13, 5, -2, 11, 24, 3, -8, -24, -8, 1, 4, -11, 4, -18, 4, 8, -7, -19, 11, 6, 4, -25, -2, 6, -19, 29, -5, 9, 24, 31, -13, -28, 7, 14, 1, 3, -22, -22, -22, -8, 8, 5, 3, 4, 8, 13, -12, -30, 9, -21, -5, 2, 21, 4, -4, 6, -14, 36, -11, 19, -8, 14, -29, -9, 2, 29, 3, -19, -39, 36, 8, -21, -13, -41, -5, -28, -2, 6, -4, -78, 28, -11, -22, -24, 2, -12, -34, 27, -2, 4, 3, 9, 3, -20, -4, 8, -26, 32, -18, 19, -11, 13, 7, 5, 5, -11, 24, -22, -2, 21, -13, 12, 16, -27, 34, 16, -4, 17, 21, 5, 5, 21, -7, 2, 4, 4, -7, -20, 12, -16, -30, -18, -9, 9, -14, -3, -2, 20, -4, 15, -18, 34, 20, 36, 14, 20, 13, 5, -19, 36, 12, 4, -18, -9, -11, 31, -28, 24, -34, -13, 1, 9, 30, -16, 29, 13, -5, -16, -30, 20, 21, 21, -10, 37, 30, 29, -21, 17, -4, -22, -4, 34, 5, -11, -20, 12, 12, 25, 0, 22, -4, -19, 2, 25, 12, -32, -39, -10, 16, -16, -6, 12, -28, -13, -4),
    (3, -53, 14, -26, -29, -1, -10, 8, 15, 18, -15, -13, -14, 17, -6, 41, 4, -11, 18, 2, -20, 14, 7, -16, 4, -8, 21, -10, -7, 22, 6, 3, -14, -12, -2, -27, -11, 24, -15, -10, -7, -1, 26, 4, -11, 1, -22, 15, 3, 2, 58, -12, -34, 17, 11, 36, -23, -24, 28, 18, 12, -41, 36, 29, -12, 1, 24, -25, -18, 0, -13, -20, 1, -12, 25, 12, -27, -4, -22, -12, -13, 1, 4, -9, -29, -13, 6, 24, -25, 4, 12, 1, 17, -25, 16, 7, 4, -14, -6, 4, -8, -4, 12, 3, -10, 12, -11, -21, 12, 27, -9, 19, 35, -8, 30, 4, -10, -7, 4, 20, 8, 7, -11, 14, -9, 10, 20, 12, -13, 12, -20, -4, 26, 9, 35, -5, -5, -4, 12, -2, 4, 0, 6, 20, 20, 17, 34, 12, -12, 19, 13, 38, 5, 15, -1, 28, -9, -15, 29, -8, -16, 8, 4, -22, -1, -18, 29, -7, -1, -16, 19, -7, -6, 9, 0, -6, -3, 6, 13, 6, -4, 14, 3, 27, -4, 23, 4, 1, -15, -12, 28, -17, -22, -18, -29, 1, -4, -14, 9, -7, 7, -1, -22, 13, -5, 14, -5, 9, -6, 27, -9, -1, -18, -25, 6, 18, 12, 6, 6, -5, -5, -16, 12, -15, -31, 1, 3, -19, 23, 10, 22, 13, 12, -12, 7, 14, -20, 3, -14, 12, 23, 14, 3, -4, 15, 38, 16, 12, 26, 18, -6, 9, 1, -15, -19, -18, -38, 16, 3, -14, -10, 0, 21, 8, 8, -6, 3, 17, -25, 7, -32, -3, 5, 27, 0, 17, -18, 11, -8, -7, -12, 7, -32, -1, 4, -20, 24, -12, 23),
    (3, -8, -10, -21, -33, -13, 8, 15, 10, -15, 0, -12, -45, -4, -13, -11, 11, -21, 21, -40, 19, 10, -31, -2, 3, -41, -11, 4, 4, 20, -27, -12, 18, 4, -21, -4, -34, -61, 30, -29, 7, 30, -26, -29, -4, -18, 19, -1, 9, -23, 23, 3, 5, -16, -33, -11, -6, -5, -12, -43, -16, 43, -49, -11, 7, -1, -2, 5, 6, 24, 13, 8, -2, -8, -13, -13, 16, 8, -14, -7, 17, -20, 8, 4, -18, -17, -3, 6, -4, -4, 16, 24, -1, 13, 0, -14, -3, -15, 26, -29, -12, -4, -5, 26, -3, -15, 5, -13, 15, 18, -9, -11, 1, -4, 3, -24, -6, -22, 13, 22, 19, -9, -8, -1, 29, 4, -13, -2, 2, -25, 24, -15, -24, -11, 10, 12, 0, -13, -34, -18, -7, 17, 29, 8, -3, -24, -6, -6, 18, -44, 23, -10, 27, 3, -5, -4, -25, 8, -7, -14, 11, -3, 14, -4, 11, -8, 33, 2, 4, -5, -17, -3, 21, -13, 20, 21, -6, -29, -17, 20, 4, -22, -30, -26, 22, 18, 4, -4, -8, -4, -3, -2, -1, -5, 15, -5, 10, 13, 3, 19, -19, -25, -6, -4, -28, 0, -24, -6, 17, 1, -11, 7, -8, -17, -11, 2, 10, 0, -2, 11, 2, -4, 17, -19, -16, -5, 39, -29, 12, 7, -26, 18, -8, -56, 13, -7, -13, 29, -24, -17, 3, 20, 12, -21, -16, 25, 0, 19, 20, 1, 17, 20, 18, -2, -5, 2, 2, -10, -4, -21, -13, -22, -33, 9, -9, -23, -4, 7, 6, -2, -5, -18, 18, -25, 27, 5, -3, -6, -1, 0, -28, -17, 3, 19, 19, 16, 3, -3, 23),
    (-11, 29, -14, 27, -16, 1, 8, -12, -17, 11, 3, 17, -15, 5, 13, 16, 12, 10, -12, 12, 8, -4, -1, -4, -13, 12, -9, 7, -3, -18, 21, 14, 16, 26, -14, 49, -7, -12, 10, -22, -25, 14, -11, 18, 9, -5, 8, -6, 30, 12, -18, -2, 20, 4, -12, -5, -25, -17, -13, -5, 4, -3, 20, 22, 9, 11, -13, -4, -9, -6, 20, -11, -5, -2, -2, 2, 7, 8, -19, 4, 22, 15, 3, 1, 5, 28, 3, -7, -7, -9, -7, 12, -10, 14, 19, 12, -3, 22, 19, 15, -20, -18, -3, -20, 2, 41, -5, 47, -12, -8, 5, 17, 8, -10, -6, 7, -12, 5, -18, -35, -32, 25, 14, -13, -1, -5, 11, 20, 9, 1, 17, 36, -28, 8, 9, -13, -3, 30, -9, 52, -1, -20, -3, 0, 15, -11, -30, 3, 3, -4, -36, -24, -8, 6, -4, -16, 6, 12, 11, 28, 14, -4, 29, 8, 11, 0, 4, -13, 1, 14, -14, 9, 6, -4, -20, -5, 13, -2, -12, 30, -23, 6, -7, -20, -2, 8, -2, -8, -7, -1, 5, -1, -11, 17, 5, 11, -20, 4, 45, -8, -13, 25, 5, -4, -3, -13, 1, 24, 5, -19, -17, -10, -21, -3, -14, -15, -22, -9, -7, -27, 22, -22, -4, 20, 20, 9, -6, 21, -7, -24, 27, -23, 0, 48, -13, 2, 10, 21, 4, 3, -10, -24, -23, -2, -16, -9, -16, -4, -10, 1, 12, -24, -21, -18, 14, 19, 12, 25, 11, 10, 8, -4, 4, -42, -2, -6, 5, -8, 7, -11, 3, 2, 22, -2, -4, 16, 5, -8, 8, 13, -27, -15, 16, -8, 6, 4, -11, 6, -5),
    (2, -22, -12, -9, -8, 15, -4, -7, 25, -12, 9, -38, -27, 2, 5, -9, -12, -14, 10, -8, 2, 7, -20, 1, -11, 11, 41, -5, -1, -1, -10, -32, 11, -16, -29, -5, 15, -3, 0, 10, 24, -8, 34, -62, -14, 32, -20, 2, -27, -5, -4, 3, 13, -21, -27, -25, 20, 14, 7, -4, 14, 5, -29, -50, -4, 17, 6, -4, 8, -3, -2, -33, 18, 7, 11, -42, -1, 14, -11, 8, -4, -4, -14, -17, 9, -20, 16, 7, 21, 5, 9, -2, -3, 11, -14, -20, -7, -20, 15, 13, 22, -5, 15, 2, -7, -21, 2, -7, -4, 10, 17, 15, -3, 6, -1, 1, 1, 4, -16, 36, -2, 13, -12, 2, 20, -4, -18, -4, 9, 32, 3, 5, -6, -5, 48, 35, 13, -28, -5, -19, -15, 25, 4, 6, -5, 28, -14, -27, 9, 16, 1, -17, 19, 7, -5, -4, -27, -2, -8, -22, 11, 20, -2, -2, -1, -3, 18, 12, 12, -8, 12, 8, -5, 18, -10, 31, -5, 20, -12, -17, -8, 13, 4, 30, -17, -8, 1, -9, -4, 1, -20, -28, -1, 8, -10, -13, -13, -14, 7, 1, -20, 2, -26, 9, -9, 7, 3, -10, -4, -20, -7, 21, -4, 1, -3, 3, -8, -4, 0, -10, -8, -1, 49, 4, -20, 18, 4, -4, 1, 14, -5, 23, -17, -32, -2, 20, -6, -31, 15, 11, 14, -17, -13, 25, 4, 3, -14, -15, 18, 28, 12, -11, -26, 3, 18, 23, 23, -7, 2, 20, 7, 8, 10, -33, 2, -16, 0, 14, 30, 13, -3, 2, 17, -19, 6, -11, -4, 6, 11, -32, 16, 17, 23, -5, 2, -5, 24, 2, -11),
    (-27, -28, -7, -8, 20, -9, -3, -19, 31, 12, -6, -3, -3, -11, -13, 14, -27, 14, 23, -15, -2, 19, -20, -20, 3, 14, 5, -19, -3, 20, -16, -3, -13, -9, -33, 14, 4, -7, -20, -26, 8, 16, -27, 28, -14, -18, -11, 0, -7, -14, -8, -8, -26, 3, -20, 3, -20, -3, -17, -18, 11, 33, 3, 20, -5, 7, -16, -1, -11, 25, -14, -12, -45, -8, -8, 36, 6, 11, -24, -18, 18, -8, 4, -4, -24, 18, -7, -16, -7, -5, -9, -16, 2, 3, 12, 17, 4, -5, -25, 3, 11, 9, 16, -25, 23, 14, 9, -7, -14, -21, -10, 23, -10, 28, 3, -14, -11, 20, -18, -7, -4, 2, -13, -4, 0, 11, -11, -7, 2, 9, -4, 8, -20, -15, -5, -30, 14, 21, -6, 19, -3, -7, -13, 11, -12, 22, -3, -2, -25, 16, -22, -34, -19, 12, 8, -6, 28, 23, -13, -2, -12, 0, 3, -2, -2, 2, -14, -49, -36, -2, -7, 26, 12, 4, -14, -20, -4, -2, -27, -17, -24, 25, 5, -13, 1, 4, 11, 3, 16, 8, -10, -3, 17, -7, 3, 4, 10, -3, -14, -6, 30, 13, 2, -18, -22, -26, -12, 0, -24, 23, 5, -15, -3, -1, -3, 4, -3, 3, -12, -20, -13, 6, 4, -12, 16, -2, 10, 21, -21, 2, 7, -11, 12, 24, 12, 11, -2, 7, -22, 2, -10, 27, -5, -11, -4, -3, -31, 3, 2, 3, -13, -21, 8, 13, 3, -11, 19, 3, 6, 4, -10, -8, 12, -23, 11, 16, -3, -2, 19, -5, -19, -7, -10, 9, -1, -8, -39, -10, 17, 7, -9, 6, -4, -17, 20, 5, 8, 1, -11),
    (6, -9, 0, 25, -18, 10, 3, 6, -7, 0, 4, 15, 5, -5, -3, 9, 5, -5, -45, 0, 9, -1, -29, -12, 6, -11, 4, 20, -26, -14, -23, 22, -1, -9, 17, 18, -13, -2, 3, 6, 0, -12, -14, 27, -11, 18, 3, 8, -7, -13, 4, 19, 8, -16, -15, -21, 27, -3, 4, 4, -8, 12, 1, 23, -11, -11, 4, 20, -2, 5, -5, 18, -2, -11, -6, 5, -5, 6, 3, 7, 6, -13, -8, 12, 12, -11, 17, -18, 9, -1, -6, -3, 5, 9, -9, -14, 19, -27, 10, 18, -21, -14, 1, -19, 28, 27, -20, -2, 28, -18, 10, -3, -23, -31, 28, -11, -12, -21, -22, 8, 11, -20, 20, 5, -25, 21, -40, 34, 14, -33, 26, 21, 11, 16, -3, -20, 20, 15, -10, -23, 20, -28, 2, -6, -28, -42, 33, 7, -14, 0, -11, 18, 23, -16, 3, 2, 45, 30, -28, -15, 24, 9, 20, 26, 4, 4, -33, -29, -7, 2, -11, -16, 11, -29, 4, -2, -1, -20, -6, 8, 5, -9, 14, -3, -13, -5, -22, 25, 28, 18, -4, -26, 8, -17, 8, -15, -1, 7, 10, -3, 2, -25, -18, -2, -7, -8, -13, -20, -14, -32, 0, -1, -18, 3, -7, 3, 2, -44, 14, 10, 17, 12, -9, -44, -9, -10, 21, -8, 19, 29, 21, 29, -15, -31, 2, -39, 15, -10, -15, 9, 0, -3, 7, 7, -20, -18, 20, 14, 11, -6, -3, 11, 13, -27, -30, -29, 7, -1, 10, -29, 14, 20, 5, 6, -9, -6, -10, -11, -2, -3, -14, -13, 5, -17, -1, 10, -20, -3, 4, 14, -17, 13, 4, -6, 15, -30, 12, -21, 17),
    (-20, 12, 3, -2, -48, -4, 12, 2, 4, 20, 17, 7, 7, -14, -39, -1, 21, 3, 18, 13, 4, 1, 8, -16, 4, 2, -19, 10, -12, 4, 15, 6, -14, -5, -10, -21, 7, -17, -3, -27, 0, 21, -17, 12, -11, -21, -39, -4, 5, 23, 38, 10, -9, 9, -4, 6, 11, 0, 25, -12, 25, 16, 3, -1, -4, 12, -14, -17, -6, -15, 15, -5, -6, 7, -21, -3, -1, -1, -15, -5, 11, 1, 31, 8, -4, 17, -11, -4, 18, 3, 5, -34, -11, 20, 10, -11, 1, -1, -13, -22, 14, 5, -16, 4, 43, -5, -9, 1, 12, 8, 5, 25, -6, -30, 34, -2, -5, 18, -19, -4, 2, 25, 3, -11, -18, -8, -16, -20, -4, 15, -1, -20, 18, -6, -37, -23, 18, -10, -12, -20, -7, -2, 4, 22, 1, -19, 35, 18, 17, 12, -9, 18, -9, 18, -12, -3, 25, 3, -27, -25, -9, -2, -1, -16, -4, -29, -25, -24, 18, -18, -24, 13, -14, 6, -14, 28, -10, 9, 25, -2, -12, 5, 16, 12, 10, 6, -21, 16, 15, 15, -4, -14, 3, 6, -5, -4, 2, 6, -5, 16, 17, -11, -2, 5, -29, -9, -20, 7, 4, 9, 1, 9, -18, 28, -23, 22, -4, -42, -12, -6, 24, 27, 3, -19, 5, 16, -17, 9, 2, 7, -5, -2, 23, 4, 16, -10, -1, -11, 4, 2, -3, 13, 9, 4, -3, 24, 0, 23, 16, -2, -3, -2, 36, -8, -23, -12, 4, 1, -2, -1, 5, 11, -3, 16, 19, -10, 16, 10, -19, 12, -10, 8, -4, -4, 7, -3, 6, 9, 20, 30, 26, -10, -8, -4, 2, -13, 4, -1, 4),
    (-27, 36, -32, 7, -1, 5, 22, 0, -6, -5, -5, -3, 1, -1, -22, -10, 0, 5, -2, 6, 18, -27, 18, -3, 2, -7, -1, -12, 9, -9, -30, -35, -12, 36, -15, 8, 1, -17, 40, -3, -5, 2, -3, 6, -33, -14, -7, 0, 1, 6, -19, 49, 10, -8, 13, 11, 21, -13, 19, -4, 6, 10, -15, -42, -21, 38, -30, -7, -23, -11, -13, -7, -9, -13, 4, -10, -18, 4, -15, -26, -7, 11, -5, 25, 17, 30, -17, 5, 10, -3, 5, -9, -10, -9, 8, 1, -5, 14, 10, 13, 5, 3, -6, 18, -13, -22, -4, 11, -26, 13, 7, -13, 21, -12, 4, -2, 13, -27, 1, -8, 22, 4, 2, -1, 5, 12, -29, 5, 10, 17, -4, 6, 34, -5, 45, 22, -4, -7, -31, -13, -16, -4, 1, -13, -10, -5, -22, 27, 20, -17, 17, -13, 36, 46, 0, -37, -15, 30, -21, -3, 3, 38, -26, 10, 33, -9, 13, -5, -21, 2, -29, 14, -4, -21, 1, 4, -8, -28, -22, 37, 11, 3, 0, -28, 21, 14, -15, -9, 0, 8, -6, -15, -1, -9, -12, 1, 4, -14, -17, 5, -6, -16, -11, -4, -2, -15, 0, -16, 9, -19, 39, -32, 5, -9, 3, 12, -14, -35, -6, 3, 21, 20, -19, -1, 20, -4, 9, 4, -12, 1, -12, 4, -1, 4, -13, -15, -8, 0, 4, -12, 11, -16, 5, -30, 4, 15, 12, 9, -7, -11, -19, -4, 20, 7, -6, -14, 33, 3, -2, -11, 2, -1, -13, -4, 17, 0, -2, -15, 8, 19, -3, -7, 10, 2, -13, -9, -3, 9, 2, 7, -17, -2, -4, 1, 9, 19, -20, -32, -8),
    (20, -22, -5, -3, 8, -20, 6, 13, 28, 2, 17, 20, -6, 19, 1, -1, 3, -1, -6, -16, -3, -22, -6, 12, 16, -8, -23, 4, -3, -13, -9, 11, 0, -19, -11, -5, -23, -4, 8, 18, 19, 14, 20, 29, -9, 24, -8, 5, 20, 9, 4, -39, 4, 6, 4, -18, 4, 4, 5, 21, -24, -25, -6, 29, 3, -4, -4, 12, -15, -12, -14, 15, 13, 12, 10, 4, 13, 34, -15, 13, 8, 4, -2, -5, 15, 4, -8, 29, 10, 8, 6, -10, 15, -23, -45, -7, -7, -45, 4, -18, -17, -4, 8, 18, 26, -4, -8, -5, -16, 17, -7, 0, 14, -18, -35, 22, 13, 3, -31, -32, 30, 4, 11, 19, -12, -12, -12, 13, -8, -43, -11, -13, -16, 27, -30, 14, 28, -1, -4, -21, -13, 37, -12, 25, -16, -28, -30, 6, 8, 19, -33, -55, 21, 28, 31, -1, -20, -19, -21, -5, -11, -3, -35, -18, -4, 10, -24, -4, 5, -4, -1, -18, -6, 10, 9, 15, -9, -19, 9, -20, 5, 10, 21, 1, 8, -7, 12, 0, 8, 10, 0, -15, -23, -3, -12, 5, -11, -1, -3, 4, 0, -29, -7, 11, -21, -2, -4, 12, 4, 4, 11, 19, -19, 14, -18, -14, 16, 2, 3, 4, 18, 4, -11, 20, -3, 9, -3, 6, -6, 7, -7, -12, 21, -5, -28, 14, -46, -4, -20, 3, 12, 9, 17, 18, -15, 37, -12, 4, 14, -15, -10, -13, 15, 0, -9, -8, 6, -7, 11, 5, -8, 1, 30, -39, 10, -13, -13, -7, -13, 3, -6, -3, 17, -4, -12, 30, -12, 13, 6, 19, 3, -26, 1, 14, 9, -13, 21, 0, -8),
    (12, -14, 6, -19, 5, -5, -1, -13, 14, 12, -29, -23, 6, 3, -9, 12, -10, 13, -21, 25, -4, 21, -7, -9, -4, 11, -4, -6, 9, -12, 14, 1, 4, -10, 5, -27, -20, -27, -15, -19, 25, 9, -12, -27, -14, -10, -6, 27, -40, 14, 16, 1, -23, 5, -11, 23, -11, 12, -21, 1, 20, -6, 21, 2, 5, 5, 9, -22, -9, -9, -16, -2, 16, -1, -15, 0, -5, 5, -9, -13, -27, 15, 9, -11, -22, -4, -15, 16, 0, -8, -5, 6, 12, 31, 22, -2, 0, 20, -4, 20, 12, -4, -4, -4, -29, -3, 18, 24, -2, -12, -8, -12, -16, 28, -4, -25, -13, -5, 28, -4, -9, -17, -8, 3, 6, 20, 28, 8, 20, 45, -1, 39, -6, 8, 12, 14, -20, -9, 33, 14, 19, -11, 1, -5, 4, 36, 3, -17, -11, 14, 40, 21, -29, -3, -3, 4, -2, 4, 13, -2, 8, 36, 28, 31, -16, 15, 4, -6, -20, 1, 24, 17, 5, -8, -3, 12, -4, 39, -21, -11, 5, 5, -3, -5, -24, 4, -10, -8, 2, -11, 5, -22, -37, 11, 22, -11, 6, 5, 25, -8, -24, 1, 5, -5, -5, -10, -36, 11, 7, -14, 6, -6, 4, -1, 6, 1, -5, -15, 17, -24, -6, -21, -9, -7, -32, 13, -3, 9, 10, 15, 17, -15, -31, 20, -6, 10, -10, -21, -11, -4, -9, -36, 9, 22, 3, -23, 26, 3, -15, -16, -6, -4, 0, -23, 8, 5, -23, 11, 13, 6, -4, 3, 2, -29, -5, -12, -11, -25, -16, -10, -6, 6, 26, -7, 9, 0, -6, -13, -11, 8, -12, 1, 6, 2, 3, -22, 27, 2, -2),
    (17, 10, 10, -6, -5, 31, -18, 15, -31, -8, 34, -4, 12, 8, -5, -39, 4, -10, -8, -31, -15, -22, 4, 5, 13, -10, 0, 6, 15, 3, 18, -4, 4, 7, 3, 6, -10, 4, 15, 33, -35, -40, 36, 4, 10, 13, 12, -30, 14, 6, -9, -28, 1, 2, 12, -5, 17, 12, 10, 4, -28, 20, 12, 22, -4, -6, 1, -9, 17, -4, 26, 19, -4, -2, 20, 4, -9, 19, 8, -25, 6, -5, -20, 10, 10, 2, 9, -6, 15, 7, 30, 13, -3, 4, 0, 3, -13, -3, 3, -16, 18, 14, -13, 8, -37, 3, -37, -4, -2, 11, 12, -5, 14, -6, -7, -13, 3, 6, 10, -13, 0, 0, -2, 25, -2, 9, 5, -1, 2, 25, 3, -6, 13, -9, 8, -2, -32, 6, 6, -26, -6, 12, 17, -20, 1, 8, -20, -28, 22, -27, -4, 14, -5, 10, -3, 5, -20, -3, 20, -13, 20, -12, 5, -7, 12, -23, -4, -2, -19, 10, 11, 13, -4, 21, 14, -34, -18, 6, -9, -23, 10, -8, -4, -28, -5, 6, -9, -34, 2, 3, 12, 11, -8, 13, -26, -6, -2, 0, 27, -7, -21, -5, -15, -11, -26, 12, 4, 4, 2, 2, 5, 0, -11, -7, 0, -7, 3, 3, 3, -7, -19, -1, 4, -11, -13, 8, 3, 24, -9, -1, 5, -1, -25, 4, 6, -17, 34, -24, 11, -6, 10, -18, -8, -23, -19, -17, 25, 16, 6, -13, -5, 10, -17, 23, 2, 2, -13, 27, 24, 24, 7, 11, 6, 7, -21, -3, 5, -15, 20, -17, 8, -15, 14, -11, 0, -10, 23, -13, 10, -8, -8, -1, 15, -1, 19, -7, 17, 26, -11),
    (-15, 0, 2, -11, 5, -32, -21, 22, -28, -6, 3, 12, -9, 22, -2, -13, 7, -4, 30, 6, -12, -15, 23, 2, -5, -20, 3, -11, -6, -5, 3, 11, -16, 11, -21, -7, -19, -22, -3, -6, -11, -6, 4, -2, 12, -3, -12, -28, 20, -14, 46, 5, -13, 6, 28, 23, -7, -3, 16, -3, -10, -5, 11, 12, -16, 10, 12, 23, 4, -22, 4, 19, -6, -4, 16, 6, 5, -6, -5, -1, 19, -29, -3, -2, -3, 11, 10, -1, 7, 6, 15, -23, -44, -2, 14, 18, -32, 30, -13, 11, 2, -16, -9, 13, -10, -14, 1, 18, 7, 9, -20, -5, 20, 35, 9, 17, -19, -14, 23, 13, -11, -14, -11, 18, -4, -11, 14, 10, -31, 19, -13, 9, 11, 2, 21, 28, -10, -6, -19, 20, -2, 20, -9, -8, 11, 5, 9, 7, 2, 4, 35, 12, 30, 18, 13, 23, -15, 3, -22, 9, -17, -2, -21, 1, 17, -4, 16, 37, -5, 11, -15, 22, -7, 12, -16, 14, 5, 5, 6, 13, 6, 6, -34, 12, 30, 19, 0, -4, -11, 15, 5, 12, -21, 4, -9, -8, -18, 8, 34, 13, -35, 5, -4, 16, -7, 1, -11, 1, -18, 0, -2, 15, -3, 15, -6, 3, 0, 8, 0, 20, -9, 1, -19, 13, -25, -10, -2, -4, -3, -1, 27, 10, -18, -18, -4, 12, -8, 18, 5, 12, 5, -20, -7, -9, -21, -7, 0, -3, 21, 7, 28, 11, 3, 11, 9, 8, -23, 4, -4, 10, -7, -1, -5, -1, -4, -17, -16, -23, -10, -8, -10, 8, 4, -13, -24, 1, -12, -2, -13, -11, 25, 3, -5, -12, 20, 8, -1, -16, 18),
    (-13, -31, 3, 16, -14, -27, 2, -8, -1, 11, 6, 28, -26, -21, -9, -3, 11, 7, -30, -13, -7, -18, -19, -16, -5, -33, -14, 2, 7, -22, -12, 23, -13, -13, -11, 7, -33, -22, -4, -8, 15, 12, -1, 29, -1, -8, -27, 26, 23, 10, -2, -2, -26, -19, -25, -21, -22, -8, 3, -12, 13, 1, -21, 15, -10, -7, 14, 9, -2, -4, -4, -14, 16, 24, -9, 17, 2, -3, -7, 7, 25, 3, 12, -1, -12, 6, -14, -8, -7, -9, 25, 18, -15, 0, 6, 6, -4, -23, 5, 10, -27, -28, -11, -13, 2, 10, -9, 26, -20, -21, -7, 13, -5, -10, -18, 25, -2, -18, -20, -33, -1, -20, -46, -10, -10, 28, 10, 28, -19, 31, -20, 8, -21, -11, -3, -13, 18, 25, -23, 61, -13, -1, -12, 20, 20, 1, -3, 37, -1, 1, -34, -12, -4, -4, -8, -36, 0, 22, -19, 33, -20, 15, 15, 11, 11, -9, 1, -5, 25, 17, -30, 26, -7, -7, -7, 2, 21, -10, -11, 28, -5, 27, 1, 7, -4, 2, -22, 51, -15, 7, -15, 12, -5, -1, 2, 0, -12, -21, 12, -13, 10, 16, 0, -22, 4, -4, -3, 12, -16, -25, 12, 7, -18, -11, -8, 1, -13, -31, 11, 1, 23, 21, -20, 10, -3, -13, 2, 12, -4, -10, -23, -28, 6, 5, -4, -14, 15, -29, 11, 3, -8, -17, 5, 0, -14, -7, -22, 9, -2, -32, 3, -1, 6, 23, -8, 0, 6, 19, 23, 5, 11, 8, 10, 3, 27, -6, -6, -9, 6, 7, 2, 3, 13, -11, 12, -11, -7, 4, 15, 22, -20, 9, 2, 29, -17, 17, 3, 2, 20),
    (-3, 3, -8, 37, -13, -14, 13, -4, -17, 14, -13, 5, -13, 26, 4, -2, 16, 5, -20, -7, -3, -8, 17, -20, 11, -20, -19, -19, 2, 27, 6, 11, 18, 13, -2, 11, 18, -13, 5, 4, -4, 15, -10, 4, 12, 30, -21, 3, -4, 21, -42, -2, -20, 1, 21, -21, -3, 23, -3, -15, 5, -14, -1, -1, -6, 19, -5, -33, 25, 23, 7, -10, 11, -18, -24, -6, 21, 18, -13, 27, -14, -14, 0, -2, -20, 5, -12, 5, 12, 7, 7, -2, -9, 6, -9, -18, 8, 17, 7, 14, -1, -16, 27, -13, 10, 23, -21, 5, -25, 18, 4, 11, 12, -2, -25, -37, 12, -8, -32, -4, 22, -10, -22, -6, -17, 25, -22, 11, 4, 37, -2, 29, 11, -12, -7, -10, 9, 43, -23, 16, 4, 3, -4, 12, -20, 3, -39, -30, 13, -17, -7, -21, -5, -9, -20, -29, -9, 27, -17, 9, -10, -28, -8, 25, -18, -12, 4, 10, 26, -1, -10, 1, -14, 25, 5, 1, -2, 18, -5, -23, -20, -28, 16, -31, -6, -5, -27, -11, 11, 21, 13, 2, -17, -1, -22, -11, -10, -34, 6, -36, -10, 18, -10, 6, -14, -14, -12, -15, -14, -13, 14, -9, 5, 7, -9, 21, -40, -19, -31, -14, 16, -2, -11, 35, 9, -1, 13, -1, 2, 4, 27, 10, 0, -26, 11, -19, -8, -27, -12, -30, 5, -17, 34, -8, -16, -6, 3, 36, -21, -57, 5, -9, 44, -7, -12, -1, -20, -13, -13, -25, 1, 33, 20, -6, -1, -8, 1, -30, -10, -9, -3, -20, 22, -8, 13, 9, -2, 18, 20, -5, 28, -11, -37, 5, 3, -37, -11, -15, -6),
    (-12, 9, 3, -10, -9, 23, -5, 12, -8, -7, 25, -7, 11, -2, 33, -23, 17, -2, -23, -18, 8, 3, 28, 7, -14, 7, -13, 5, 5, -20, 27, 16, 23, -17, 21, 2, 10, 8, 2, 12, -17, -27, 16, -41, 4, 32, 26, -29, -6, -12, -21, -20, 24, -34, 9, 7, 3, 8, 12, -7, -11, -16, 6, -15, 19, 11, -2, -6, -5, -14, -7, 0, -5, -10, 28, -24, 7, 30, 9, -10, -3, -18, -7, 5, 22, -3, -6, -15, 2, 0, 9, -12, -12, -2, -8, -17, 12, -14, 16, -22, 2, 31, -36, 33, -3, -24, 5, -4, 5, 10, 9, -25, 5, 12, 10, 2, 1, -15, 18, 1, -5, 13, 19, 11, -10, -22, 42, 8, 10, -26, -2, 13, -13, 27, -6, 9, -20, 2, 19, -13, -2, 29, 27, -5, -8, -3, -15, 4, 15, -23, 23, -35, -12, 9, 7, -20, -5, -24, -13, -18, 20, 6, -21, 11, 7, -4, -4, -42, -7, 21, -4, 4, 25, 1, 19, 0, 13, -25, 0, -10, -1, -4, -17, 7, -9, 0, -1, -36, 8, -10, 1, -8, -4, -8, 16, -13, 10, 26, -6, 1, 18, 4, -4, 1, -24, 20, -20, -11, -19, 8, 2, -11, -4, 28, 1, -12, 13, 20, 13, -14, -3, -11, 8, 5, -20, 0, 4, 7, 11, -24, 3, -13, -2, 18, 2, 6, 15, -20, 19, 15, 27, -8, 0, 12, 20, 0, -12, -11, -11, 12, -11, -27, 2, -1, 5, -17, -10, 8, -16, -3, -2, -3, 6, -41, -18, 33, -20, 32, 12, 10, 4, -8, 0, 12, -4, 13, -8, 26, -12, 21, -9, 9, -8, -5, -17, -2, 5, -2, -16),
    (10, 10, -6, 3, 5, 11, 5, -12, 6, 16, -25, -4, 5, -18, 10, 2, -16, -44, 9, 23, -4, -4, -10, -17, 0, -2, 18, -21, -12, 15, -21, -11, 0, -5, -28, 4, -7, -32, 12, -20, -4, 0, -17, 26, 18, -27, 1, -4, -9, -51, 13, 17, 7, 3, -14, -19, -9, -1, 4, -6, 15, 35, -23, -6, 9, 20, -31, 10, 10, -16, -13, -2, -8, -4, 1, -7, 7, 0, -10, -18, 11, -57, 4, 20, 11, -5, -31, 22, 39, -25, 11, 14, 14, 36, -9, -11, 21, -20, 21, -44, 2, -2, 6, -17, 2, 5, -19, -26, 0, 12, 7, -4, -34, -11, 13, 10, -3, 2, 26, -8, 7, 17, 10, -7, 23, -2, -6, -37, 12, 8, 17, -24, 12, -8, -17, -26, -14, -3, -26, -31, 16, -11, 12, 2, -37, -14, -11, 12, -18, 7, 4, -5, -5, 24, 2, -4, 20, 10, 15, -36, 4, 4, -23, -28, 36, -11, -13, -20, -14, 9, -22, -7, 13, -10, 15, -1, 5, -9, 3, 23, -22, 4, -16, -10, -9, 0, 14, 7, -10, -1, 7, 9, 8, 13, 18, -1, -7, -4, -15, 5, -1, -12, 29, 0, -9, 16, 19, 9, -9, 12, -1, -7, 12, 29, 11, 11, -9, 7, 7, -18, -13, 13, -11, -5, 5, 13, 20, -16, -4, 12, -32, 4, 11, 4, 33, -12, 17, 12, -1, -12, -3, 21, -14, -7, 12, 19, 19, 11, 23, 10, 20, -4, -3, 8, -16, -14, 8, 11, -6, -5, 13, 1, 8, 24, -9, 9, 27, 19, 4, 8, -3, -16, -4, -4, -1, -18, -2, 13, 4, 11, -12, 28, -3, -13, 23, 17, -8, 19, 9),
    (6, -3, 12, -24, -3, 2, 4, 20, -3, -13, -10, -15, -8, 5, 11, 26, -23, -19, 0, -8, 9, -11, 1, -10, 19, -9, 17, -14, 6, 3, -19, -30, 0, -21, 16, -45, -5, -5, -4, -3, -10, 0, -43, -17, 20, 24, 20, 7, -50, -4, -24, 11, 3, 4, 6, -28, 19, 17, 10, -15, 13, 16, -3, -20, 6, 13, -14, -13, 7, 2, -15, -2, -26, -14, -36, 36, 39, 12, 21, -14, -20, -3, -9, 5, -15, -10, -3, 17, 6, 16, 2, 0, 7, 11, -5, 0, 26, 17, 24, -21, 6, 8, 3, 15, 5, -14, -10, -45, 1, -2, 26, 12, -8, 3, -18, 5, 3, 18, 18, 9, 2, 9, 9, 5, -13, -3, -5, -23, 8, 21, 30, -34, -7, 14, -34, 13, 3, -34, -4, -32, 7, 26, -8, 8, -44, 21, -4, -11, 1, 13, 11, -12, -7, 17, 22, 16, 27, -18, 11, -37, 1, -10, -30, -53, -7, -10, -29, -20, -8, -5, -4, -8, 18, 10, -2, -25, -3, 5, -5, 8, -17, -3, -20, -4, -12, 10, 5, -14, 33, 12, 4, -20, 1, 6, -13, 14, -21, 14, 2, 8, 3, -3, 11, 19, 18, -2, 6, 2, -3, 21, -11, 11, -1, -16, -13, -2, 24, 7, -6, 0, -7, 2, -13, 11, -12, 20, -2, -21, 4, 12, 7, 29, 9, -4, 9, 9, -35, 12, -28, 19, -9, 15, 12, 25, 4, 29, -9, 8, 11, -3, 5, -24, 20, -13, -14, 12, 10, 21, -4, -26, 6, -17, -9, -9, -17, -5, 10, 33, 2, 18, -24, -22, 35, 15, 25, 22, -24, 8, 2, 9, -34, -23, -22, -4, 16, -2, -4, 0, -25),
    (-10, 34, -1, 3, 5, 6, 9, -21, -4, 4, -33, -11, -16, 19, 27, -18, -5, -14, 5, -35, 13, -39, 1, 11, 1, 5, 10, -18, 14, -28, -9, -10, 17, -10, 20, 15, -6, -5, 11, -13, -6, -2, -26, -14, 20, 23, 12, -13, -4, -12, -32, -14, 18, -30, 3, -10, -1, 0, 10, -8, 4, 0, 4, -26, 35, -16, 27, 4, 9, 3, 12, 20, 2, -17, -12, -15, 16, 18, 22, -4, -10, -4, 2, 5, 15, -16, 12, 5, 10, -12, 1, -8, 7, 30, 3, -18, -7, -17, 24, 24, -10, 13, -18, 1, 8, -5, -10, -17, 3, 6, 39, -4, 4, -12, -21, -4, -9, -2, -8, -2, -15, 9, 22, -9, 15, -25, -7, -7, 23, -59, 50, 7, -2, 16, -21, 7, 23, -4, -13, -28, 25, 8, 18, -16, -25, -22, -5, 2, 21, -11, 10, 7, -8, 4, 22, 3, 22, 3, 3, -22, 6, -38, 4, -14, -7, 3, -5, 10, -11, -19, 15, -7, 5, 0, -6, -29, 5, 0, -4, 12, 2, -26, -6, -30, 0, -13, -20, -15, 18, -8, 2, -12, 9, -17, 4, 1, -1, -13, -3, 8, 33, -2, 2, 0, 27, 11, 23, -3, -6, -20, 13, 5, 11, -17, 20, -13, 0, 2, 7, 9, -4, -5, 29, 11, 15, -29, 4, -19, -1, 22, -10, 9, 36, -9, 20, -17, 14, -11, -1, -20, 15, 6, 7, 3, -4, -8, 2, 8, -9, -13, 11, -8, 17, 5, -20, -3, -7, 12, 0, 1, -5, 3, 13, -44, -29, -26, 14, -8, -6, 0, -4, -15, 24, -12, 12, 21, -29, 9, 26, -15, -25, -14, 4, -2, 28, -17, 8, 28, -14),
    (28, -31, -3, 4, -25, -1, -14, -29, 36, 24, -33, -6, 19, -21, 28, 21, -27, -38, 1, 8, -4, 24, -22, -1, -13, -1, -12, -22, -11, 27, -35, 0, 11, -44, 16, 6, -10, -12, -23, -20, 21, 16, -4, -11, 28, -10, 24, -5, -42, -52, 33, 8, -8, -18, -6, 4, -31, 1, 2, -6, 25, 18, -22, -8, 12, -2, 3, 0, 13, 2, 9, -13, 2, 8, 3, -3, 20, -20, 21, -37, -11, -21, -5, 12, -15, 9, -16, 0, -5, -5, 11, -11, -2, 9, 5, 5, 5, -21, -2, -22, -8, 11, -29, 4, 9, 10, -31, -4, 26, 15, 1, 7, 21, -4, 0, -4, -6, 3, -10, 3, 8, 5, -13, 3, 0, -9, 5, -7, -3, -27, -7, -39, -3, -13, -20, -15, 10, -25, 0, -11, 8, 25, 13, 19, -11, -2, 36, 13, -21, 21, -5, 6, -20, -6, 14, -2, -38, -28, 34, 13, -11, 1, 17, 10, 10, 12, 3, -10, -5, 24, 1, 7, 8, -8, 0, 7, -9, -18, 0, 35, -6, 7, -19, 23, 12, 8, 13, 5, -18, 13, -2, -13, -5, 13, -3, 4, -16, 15, 8, 7, -24, 14, -14, 11, 9, 11, -20, -5, 27, -4, -9, -9, 4, -8, 2, -9, 3, -26, 10, 21, -6, -5, 25, 14, -24, 15, -6, 3, 7, 17, 10, 7, -19, 5, -2, 18, -15, 9, 3, 30, 18, 19, -7, 8, -6, 26, 1, 11, 20, -4, -11, 14, -19, -13, 17, 7, 9, 8, 16, 7, -6, 0, -25, 11, 24, -25, 3, -13, 3, -12, 7, -1, -7, -25, 2, -29, -8, -14, -34, -14, -1, 3, 9, 9, -3, 19, -1, -33, 25),
    (3, 21, -22, -19, 11, -25, 3, -31, 11, -21, -3, -17, -7, -4, -4, 9, -38, -1, -4, 8, 20, -1, -6, -7, -7, 22, 14, -29, 2, -24, -13, -22, 9, 20, -6, 1, -5, -3, -14, -33, 8, -5, -12, 17, -3, 6, -12, -16, 2, 5, 38, -28, -20, -20, 10, 0, -22, 3, -38, -19, -16, 13, 3, 2, -22, -28, -22, 33, -26, 2, 19, 9, -27, -3, -4, 20, -17, 0, -24, -30, 20, 14, 2, -18, -12, -22, -6, 13, -25, 0, -20, 26, 1, -9, -8, 3, 5, 22, 15, -4, -7, -5, -5, 13, -22, -13, 27, -3, 10, 10, -4, -43, 10, 1, 8, -9, 0, -10, 19, -12, 9, 11, 13, 7, 21, -10, -1, -1, 6, -6, 12, 4, -6, 21, 20, 36, 0, -12, 41, -12, -7, 22, -12, -20, 23, -4, -10, -8, 13, -7, 22, -7, 35, -3, 19, 12, -5, 5, -20, -2, 3, 1, 10, 9, 3, 7, 26, -4, 0, 3, 23, -23, 4, 3, -11, 3, -20, -14, -15, 1, 3, -27, -8, 27, 22, 9, 21, -12, -24, -30, -36, 13, 19, -35, 15, -9, 10, -5, -2, 13, 32, -15, -5, 1, 14, 7, -12, 14, 0, -14, -5, 9, 0, -26, -12, -13, -4, -13, -5, 5, 4, -21, 13, -19, 10, -24, -8, 3, -3, -20, -22, 12, 18, 8, -19, -11, -8, 23, -20, -12, -24, 13, -10, -21, 5, 7, -6, 1, 12, 10, -17, -16, -46, -13, -15, -27, -3, 16, -15, -24, 12, 4, -8, 19, -24, -3, -20, 32, -13, 22, -22, 7, 8, 4, 4, 1, -2, 29, -6, 7, 9, 5, -16, 41, -12, 16, 17, 16, -12),
    (-12, -12, 1, 4, -13, -1, 9, -12, -15, -3, -23, 4, -7, 7, -8, 13, -3, -12, -13, 3, 3, -15, 11, 6, 7, -9, 15, -29, -12, 27, 15, -3, -21, 12, 6, -19, 3, -11, 19, -11, 4, -13, 6, -5, -23, 0, -29, 12, 4, -3, -9, 28, 7, -13, 12, 22, 11, -15, 7, -20, -1, 4, -1, -5, -30, -7, -5, -9, -4, -2, 6, -5, 4, -22, -22, -2, -25, -13, -21, 23, -1, -4, -4, 14, -20, -17, 8, 18, 22, -16, 5, 17, -7, -17, -13, -12, 12, -2, 6, -40, 3, 12, 6, -15, 15, -10, -7, -14, 13, -30, -11, 10, -7, 21, 13, -10, 4, 12, 3, 13, 10, 0, -4, 12, 14, -4, 21, -36, 10, 29, 10, -40, -4, -2, 36, -12, 20, -26, -3, -27, -22, -12, -22, 15, -7, 16, 33, 3, 11, 0, -4, 30, 16, -16, -22, 8, 24, 12, 13, -33, -4, -12, 7, -22, -6, -14, 20, -19, 18, -21, -12, -16, -13, 1, -18, 3, 9, -3, 10, 19, -13, -9, -1, 17, 13, -4, -29, 23, 11, 12, 17, -8, 16, 5, 18, -10, 15, 0, -11, 10, -2, -33, 5, 12, -18, -4, -25, -30, -15, 7, 9, -21, -5, 1, 22, 9, -5, -4, 8, 0, 29, 1, -13, -17, 8, -3, 18, -3, 7, -3, -7, -3, -20, -46, 3, -20, 12, -29, -25, -32, 17, 4, 30, -18, -36, -6, 19, 37, 3, -14, -9, 1, 34, 15, 6, -44, 12, -1, 27, 21, -2, 11, -15, 16, -17, -37, 7, 7, -6, -10, -10, 6, 8, 11, 11, 1, -38, 11, -2, 14, 5, -7, 7, 17, 23, 5, 21, -20, 20),
    (3, -5, 15, -1, 11, 1, -3, -3, 6, -3, -29, 12, -5, 25, 14, 25, -10, 5, -8, -1, 1, -23, 1, -15, 12, 23, -3, -48, 33, 6, -26, -7, 6, -46, -9, -7, 21, -25, 5, 3, 24, 4, -36, -21, 4, 22, 2, 29, -44, -15, -6, 9, -5, -5, 18, -37, 27, 53, 24, -38, 19, 9, -30, -21, 2, 12, -4, -18, 30, 0, 15, 4, 4, 5, -25, -1, 2, 10, 8, 19, -19, -16, -36, 28, 4, 11, 2, 3, 29, 12, 10, -15, 7, 12, -2, -6, -5, -5, 0, -7, -1, -6, -16, 2, 0, -23, 11, -6, -43, 20, -24, -11, -3, 20, -1, -11, -7, 0, -15, -1, -21, -4, -5, 2, -8, -3, -16, -8, -7, 14, -4, -26, 6, 20, -53, 20, -4, -31, 12, -12, -15, 7, -13, -19, -2, 28, 13, -28, -16, -2, 12, -6, -31, -21, -3, -4, 21, 4, -23, -13, 3, -6, 10, -24, 20, -4, 15, 28, 16, 2, -6, -1, -21, 6, -1, 9, -31, 2, -11, -4, 6, -17, 6, -25, 6, 9, 6, -8, 13, 18, -19, -23, -23, 19, 5, 5, -3, -7, 9, 2, -11, -16, 11, -10, -5, -24, -3, 8, -1, 7, -6, -9, 4, 15, 1, -6, -10, -1, -5, -11, -10, 24, 10, -2, -14, 14, 11, 11, 0, -11, -17, 9, -24, -3, 21, 4, -23, -33, -13, 1, 10, 5, 7, -1, 4, 9, 7, 13, -8, -20, -19, 1, 7, 12, -29, 13, 5, 12, 7, -6, -2, 5, 10, -2, 2, 6, 8, -25, -34, -2, 1, -2, 11, 12, -7, 6, -1, 15, 21, 5, 6, -16, -6, 20, -8, 3, -11, -7, -5),
    (-22, 9, 0, -7, 4, -11, 22, 26, -20, -12, 1, -14, -4, 17, 12, -10, -25, -4, 19, 8, 12, -10, -2, 5, 34, 9, -24, -3, -4, 31, -12, 12, -19, 18, -10, -14, 18, -20, 34, 15, -22, -17, -21, -23, 12, 4, 21, -18, 9, -7, 18, 4, 22, -21, -10, 14, 46, 16, -6, -4, -20, 32, -12, -6, 6, 2, -1, 4, 47, 11, 30, 14, 0, -4, -19, -8, 6, -11, 16, 9, -5, -12, -8, 24, 21, -45, 8, -11, 28, 1, 21, 5, -17, 23, 3, -14, -9, 20, 11, -6, 2, -5, -26, 20, -15, 4, -34, -30, 0, -3, -5, 1, 0, -4, 2, -11, -21, 7, -11, 0, 14, -19, 1, 33, 12, 33, -24, -9, -15, 20, -13, -20, 13, -23, 25, 10, -13, -23, -15, -27, 11, -13, 7, -6, 5, -3, 15, -1, -7, 6, 17, 5, 30, 6, 6, 21, -10, 24, 3, -8, -6, 8, 17, -11, 29, 0, 4, 37, -18, -14, -12, -16, -4, -1, 5, -7, -1, 1, 3, 11, -10, -13, 2, -17, 18, 7, 5, 15, 20, 18, 3, -4, -28, 2, 4, -11, -15, 6, 5, 12, -25, -15, -12, 9, 18, -11, -28, 8, -5, 9, -1, 16, -19, -6, -34, 18, 3, 4, -1, -1, 2, -4, 4, -21, -45, 0, -11, -11, 1, 6, 8, -11, -11, -22, -8, 0, 15, 2, -9, -1, 13, -7, -20, 9, -30, -2, -13, 23, -12, -4, 24, 27, 1, 3, -15, -15, -6, 28, 22, 9, 3, 10, 29, 37, 3, -13, -5, 10, 15, 23, -19, 37, 10, 5, -11, 2, -17, 25, 13, 12, 5, 9, 17, 17, 4, 3, -3, -9, -4),
    (1, -2, -15, 4, 17, -10, 3, -15, 17, 20, -19, 16, 8, -40, -3, 5, -5, -21, -20, 21, -10, 19, -13, -10, 17, 4, -7, -8, 14, -1, 13, -3, 21, -20, 13, -12, -18, 10, -27, -4, 13, 12, -7, 6, 33, -16, 4, 24, 5, -21, -13, -11, 0, 4, -17, -19, -12, -12, -13, 17, 25, -31, 20, -3, 4, -23, 9, -13, -4, -13, -11, -28, 1, 13, 9, -2, 12, -2, -2, -18, -11, 1, -1, -5, -1, 10, -8, -15, -14, -2, -15, -5, 30, -4, 23, 8, 5, -43, -7, 11, -1, 18, -35, -20, 12, 2, 3, -11, -2, 4, 20, 19, 10, -25, -23, 31, -6, 9, -26, -16, -31, -11, -3, 13, -9, -12, 6, -3, 8, -33, -11, 10, -13, 22, -35, -7, 12, 13, 1, -10, 36, -4, 36, 13, -32, -10, -26, 36, -12, 30, -12, -20, -35, 11, 10, 4, 8, -33, 4, -11, 27, 6, 18, -40, 6, 15, -39, -21, 6, 17, 5, 2, 21, 10, 17, 9, -15, -1, 18, -13, 5, 9, 7, 17, -13, 10, 22, 13, 26, 4, 10, 6, -9, -5, -54, -1, 1, -2, 14, -13, 2, 17, -11, 5, -30, 36, -9, -8, 5, -5, 14, 6, -1, -19, -20, -10, -12, 6, -16, -17, 10, 1, 0, 3, -29, 4, -20, 10, -13, -14, 10, 6, 4, 7, -10, 4, -20, 29, 21, 3, -6, 3, -19, 17, 2, -1, 0, -2, 31, 12, -24, -21, -59, -10, 10, 1, 9, -13, -7, 5, -5, 20, -7, 15, 7, 3, -5, 3, 5, 23, 25, -1, 14, -8, 5, -11, -9, 1, -12, 0, 4, 8, 31, 12, -9, -12, 5, -5, -10),
    (3, -42, 6, -3, -20, 11, 3, -1, 21, 27, 2, -3, -12, 24, -17, 6, -6, -16, -24, 8, 10, 12, -10, -10, 6, -10, -1, -30, -2, 11, -21, 5, -3, 10, -9, -22, -6, 19, -29, -21, 16, -10, -16, -13, -4, 27, -4, 23, -17, -6, 1, 2, 6, 28, -8, -27, -28, 20, 10, -22, -6, -11, -9, -8, -3, 1, -9, -33, 4, 18, -25, -35, -23, 15, -29, 11, 20, -13, -12, -7, -21, -20, -3, 6, -21, 17, -16, 5, -19, 16, -2, 11, -3, 5, 0, 2, -11, 48, 3, 13, -12, 12, -28, 13, -20, 23, 18, -30, -13, -17, -8, 26, -7, -4, 10, -10, -1, -18, 10, -1, 13, -28, -15, 12, 29, 12, -18, 16, -15, 43, 5, 10, -15, 7, 15, 14, 23, 17, 16, -30, 2, 12, -12, 31, -20, 37, -20, 4, 14, 21, 5, -3, 3, 1, -12, -25, -31, 10, 0, -8, -4, 24, -1, 18, 2, 5, 1, -49, 18, 15, 3, 0, -1, 4, -16, 13, -4, 2, -16, -11, -11, 27, 7, -23, -27, 22, 2, 4, -13, 15, -7, 7, -10, -2, 3, -2, 9, -10, -9, 5, -14, 15, -16, 6, -18, -5, -7, -37, 36, -26, 0, 20, -21, -3, -1, -2, -12, -21, -2, -5, -1, -1, -23, -7, -14, -17, -5, 4, -7, -19, 9, -3, 21, -10, -21, 37, -29, -41, -11, -6, 9, -5, -10, -33, 8, -23, -13, 19, 4, -27, -28, -21, 13, 14, 5, 5, 16, -5, -9, -4, -19, -8, 0, -15, 0, 22, 4, 3, -17, 23, -16, -15, -12, 18, -12, -9, 11, -2, -22, -15, -16, -4, -17, 9, -8, -16, -16, 13, -16),
    (4, -18, 12, 12, -12, 4, -8, 28, -5, -28, -6, 13, -5, 16, 3, 7, 20, 20, -18, -35, -8, -14, 10, 2, 13, -42, -21, 9, -12, -4, 23, 6, 18, -8, -10, 12, -48, -10, 11, 21, 11, -20, 37, 5, -31, 24, -11, 4, 13, 35, -5, -48, -3, 14, 14, -29, 4, 1, -1, 18, -2, -24, 35, -4, -9, -6, -17, -14, -17, -14, 27, -9, 13, 7, -9, 6, -13, 15, -25, 2, 10, -26, 0, 15, -27, -17, -5, 17, -6, -5, 8, 0, -4, 0, -16, -14, 5, -6, 11, -3, -2, 6, 1, -21, -19, 5, 11, -11, 26, 8, 39, 5, -5, -5, -12, 4, -8, 11, 5, -7, -24, 6, 28, 19, -2, -16, 4, -14, 17, -4, 32, -27, 0, 21, -30, 21, -20, -20, 3, -22, 8, 20, 10, -20, 5, -4, -11, -12, 14, 6, 11, 6, 0, 11, 21, 20, -11, -19, 25, 13, -5, -1, 14, -19, -23, -14, 24, -7, -32, -18, 11, -23, -21, 9, 10, 10, -1, -2, 9, -18, 11, 13, 2, 21, 13, -13, -33, -11, 30, -13, -23, 23, -36, 12, -19, -19, 0, 2, 18, -5, -5, 14, -22, -5, -24, 18, -10, 12, 2, 15, 9, 7, 5, 28, -9, -4, 10, 7, -4, 0, -11, -3, 0, -2, 1, -23, 3, -14, 4, 2, -24, 5, 12, -7, -30, -10, -16, 32, -22, -5, 8, 8, -13, 3, -15, 33, 22, 12, 16, 18, 22, 10, 10, -2, 9, -17, -13, -18, -32, -13, -5, -12, 20, -21, -21, -24, -21, 8, 9, 7, 11, -29, 35, -37, 7, 17, -10, -39, 0, 16, -10, 1, -10, 8, 4, -3, 4, -20, -11),
    (-19, -33, 21, -22, -44, 20, -21, 8, 14, -24, -4, 40, -22, 26, -21, 29, 8, 23, -18, -25, -6, 31, -19, -3, -12, -21, -3, 2, -16, 2, 20, 23, -27, 3, -32, -12, -17, -16, -4, -7, 25, -29, -20, -4, -28, 20, -33, -3, 4, 10, 21, 10, -20, 2, -4, -13, -15, -17, -4, -33, 1, -5, -29, -4, -22, 9, -20, -33, 4, 3, 18, -11, 2, -2, -15, -19, -40, -12, -28, -5, -19, 9, -1, 12, -19, -16, -2, 12, -2, -15, 21, 18, 12, -25, 2, -11, -7, -24, 7, 22, -29, -1, -7, -6, -9, 11, 16, 14, -1, 2, -9, 4, -2, 6, -28, -10, -20, -4, 21, 12, -12, -21, 8, 13, 17, -15, 2, 22, -4, -3, 5, 24, -20, 5, -3, 12, -16, -14, 23, -6, -12, 36, -4, -13, 23, 40, 5, -18, -2, 1, 33, 7, -12, 0, -5, 38, -10, -21, 41, 4, -5, -4, 12, -17, 4, 4, 18, 32, -14, -21, 9, -13, 8, 32, -4, 18, -8, -6, 5, -11, -21, -4, -4, 3, -3, 4, 1, -5, -22, -30, 18, -17, 2, 4, -5, 14, 0, 5, 9, -22, -3, 27, 16, -14, 1, -4, 11, 11, -6, 3, 3, -11, -14, 3, 16, 10, 5, -2, -7, -11, 2, 4, 0, 19, -4, 9, 11, 21, 0, 2, 6, -9, -3, 40, 12, -15, -7, 10, 8, 5, -16, 9, 10, -23, 12, -5, 26, 15, -11, -11, 8, 4, 19, 4, 2, 14, 15, -4, 15, 26, -4, -28, 2, -31, 20, 26, 0, -8, -5, 10, -3, -7, 11, -2, 11, 22, -15, -13, -2, -12, 8, 11, 1, -11, 12, -24, 8, 3, -4),
    (-5, -33, 17, -21, 3, 17, -12, 20, 11, -18, 12, -23, 4, 28, 25, 9, 8, -19, -24, 0, 18, -5, -5, 3, -5, 27, 14, 12, -33, -28, -10, 1, 11, -46, -4, -43, -4, 23, -4, 24, 12, -24, 29, -20, 0, 24, 8, 4, 11, 0, -5, -4, 11, -14, -11, -3, 9, -22, 8, 31, 7, -21, -3, -8, -15, 3, -2, -24, -5, -3, -9, -20, 12, -11, 17, -17, -1, -7, -5, -24, 17, -10, 19, -9, -23, -11, 0, 12, -10, 15, -13, 30, 4, -8, -9, -3, 42, -51, 20, 11, -5, 11, -15, -4, 20, 7, -5, -21, -1, 10, 0, -2, -11, -3, -21, -19, 13, 11, -19, -17, -12, -4, -3, 1, 13, -11, 2, -19, 16, -29, -5, 2, -26, 14, -13, 12, -21, -19, 19, -15, 2, 5, 10, -57, -1, 12, 16, -47, 10, -21, -4, 4, -4, -18, -26, 6, 24, -16, 10, 4, -37, 6, 11, -4, -16, 4, 43, 1, -21, -1, -5, -13, -17, 17, -17, 12, 16, 16, 27, 12, -3, 4, 15, 17, -7, 4, 10, 1, -26, -16, -27, 4, 20, -4, 1, 2, 4, -19, -25, 17, 8, 10, 4, -24, -5, -12, -1, -12, -3, -2, -4, -8, 19, -18, -4, -12, -7, 3, -6, -1, -2, 11, -12, -27, 21, -5, 26, 9, -2, 19, -13, 5, -24, 4, 9, 13, 16, -2, 21, -35, 16, -1, -1, 3, -5, -3, 4, 9, -7, 8, -3, 10, 16, -18, 10, -11, -19, 15, 30, -11, -2, 3, 30, 20, -58, -1, 2, 3, 0, -14, -25, 19, 10, 8, 42, 14, -35, 6, 10, 21, -7, 6, -1, -6, 7, -8, 2, 36, -17),
    (10, 3, -4, -4, -13, 13, 0, 48, -29, -44, -10, -16, 1, 36, 11, -40, 32, -7, -11, 6, -4, -37, 21, 11, 14, -21, 4, 28, -24, 8, -2, 20, -17, -1, -10, 4, 19, -8, 19, 40, -35, -11, -17, -5, 6, 38, 15, -35, 25, -2, -4, 21, -3, -29, 36, -1, 10, 11, 20, 22, -21, 8, 19, 5, 1, -2, -29, 7, 11, -3, 3, 31, -12, -8, -12, -8, 19, 25, 16, 13, 3, 2, -2, 4, 11, 2, -13, -18, 4, 15, -3, -38, -12, 15, 12, 4, 9, 5, 4, -6, -10, -4, -9, 27, -28, -25, 3, 7, -5, 20, -1, -29, -5, 4, -5, -37, 5, -29, 19, -12, 6, -19, 9, 27, 5, 5, 28, 13, -12, 4, -20, -14, 8, -14, 11, 36, -21, -18, 7, 1, 4, 23, 4, -34, -2, -1, -12, -13, 3, -13, 41, -17, 18, 3, -2, 22, 5, 6, 6, 11, -21, 1, -62, -11, 9, -7, 24, 22, -13, -7, 8, 10, -21, 19, 19, -22, -1, -4, -12, 11, 13, -3, -24, 0, 0, 7, 3, -31, -1, 20, 14, 10, -1, -9, 0, -7, -9, -13, -6, 10, -10, -10, 4, 4, -1, 10, -9, 10, -15, 7, -16, 5, 12, -1, 18, -17, -1, 20, 12, 14, -2, 5, 16, 13, -11, -4, -14, -24, -1, 8, 0, 10, -17, -11, -6, 9, -17, 12, 4, 4, 11, 12, -13, 8, 0, 25, -6, -18, -4, 4, -6, -5, -2, 8, 7, -1, -19, 3, -5, -12, 0, -12, 2, -2, 3, 16, -4, 1, -27, 16, 8, -6, -5, 7, -6, 16, -10, 31, -21, -15, -6, -5, -6, -27, -2, 9, 14, 0, -6)
  );
  ----------------
  CONSTANT Flatten_1_Columns : NATURAL := 2;
  CONSTANT Flatten_1_Rows    : NATURAL := 2;
  CONSTANT Flatten_1_Values  : NATURAL := 32;
  ----------------
  CONSTANT NN_Layer_1_Activation : Activation_T := relu;
  CONSTANT NN_Layer_1_Inputs     : NATURAL := 128;
  CONSTANT NN_Layer_1_Outputs    : NATURAL := 10;
  CONSTANT NN_Layer_1_Out_Offset : INTEGER := 6;
  CONSTANT NN_Layer_1_Offset     : INTEGER := 1;
  CONSTANT NN_Layer_1 : CNN_Weights_T(0 to NN_Layer_1_Outputs-1, 0 to NN_Layer_1_Inputs) :=
  (
    (-2, 29, -35, 26, -6, -37, -45, -13, 9, 28, 6, -44, 9, -44, 20, 22, -50, -5, 6, -5, -2, 9, -33, 42, 2, 11, 42, -27, -15, -8, -28, -14, -4, 2, -1, 17, 10, -6, -27, 4, -14, 3, -17, -23, 11, 5, -8, 27, -12, 11, -9, 2, 7, -3, 11, 6, -6, -5, 2, -2, -1, -3, -26, -18, 35, -2, 17, -1, -3, -34, -24, 5, -3, 10, -8, -16, -2, -26, 14, 8, -19, -20, -10, -12, -6, 12, 19, -19, -25, -9, 4, -10, -27, -1, 7, 10, 2, 2, -8, 3, 12, -8, -22, -8, 13, -6, 3, 0, -6, 1, 8, 6, -10, 4, 4, -2, -1, 18, -25, 12, -5, -5, 4, -19, -3, 16, -2, -2, 14),
    (19, -13, 30, 6, -1, -9, 18, 24, -27, 9, 2, -10, 42, 14, -57, -18, 12, 4, 22, 18, 8, -26, 5, 12, 20, -13, -8, 18, -24, -7, 6, -14, -1, -5, -9, 11, -7, 12, 5, 11, -18, -2, -13, -15, 15, -36, 19, -11, 7, -14, 16, 24, 15, -16, 15, -2, 7, -24, -6, -10, -19, 5, 10, -6, -10, 10, 5, 3, 0, 11, -4, -17, -8, -4, 0, -12, 5, 7, 12, -3, 8, 7, 14, 7, 1, -22, 18, 10, 0, 16, 2, 14, 17, -10, -8, -20, 8, -11, 9, -14, -3, 5, -7, -4, -1, 10, -10, -7, 15, 2, -14, -10, -7, -13, -7, 9, 25, -3, 12, 4, -6, -7, -6, 9, 18, 5, -16, -9, 3),
    (20, 7, -9, -22, 6, 13, 5, 13, -17, 14, 0, 14, -21, -30, 19, -14, -10, 10, 9, 29, 30, 14, -26, -25, 27, -25, 26, 11, -9, -32, 9, -43, 19, -7, -31, -5, -18, -14, 3, -8, -12, -2, -10, -10, -3, -14, 6, -11, 6, 6, 3, 22, 29, -4, 9, -13, 6, -18, 18, -10, 2, -18, 10, -31, -11, -7, 5, 1, -5, 1, 10, 22, 12, 16, 22, 12, -2, -18, -13, -1, -14, 9, -7, 16, -10, -9, 3, -13, 22, -11, 14, 17, 4, 8, 10, -10, 0, 11, -4, 1, -4, 8, -3, 12, 3, -3, 2, 3, 2, -11, -11, -15, 5, 4, -6, -1, 1, 4, -6, -2, 3, 22, 14, 9, -12, 9, 4, -1, -21),
    (3, 10, 31, -17, -25, 43, -2, 20, 15, -17, -29, 6, 6, -5, -10, 34, 18, -39, -10, -42, -2, 17, -19, -35, -25, -47, 10, 18, 2, 26, 0, -1, 10, 15, 7, 11, 9, 16, -17, 1, 12, -5, -24, -21, 16, 21, 0, 21, 7, -20, 7, -8, -15, 14, -2, -2, 3, -20, -5, 13, -1, 20, -3, 6, -8, 2, -6, 2, 22, 6, -9, -14, -13, -20, -8, -14, -7, 1, 16, 20, 17, 0, 27, -32, 3, 24, -19, 13, -7, -10, 7, -25, -17, -26, -17, -22, 0, -4, 0, -22, -2, -3, -9, -16, 10, -11, -3, 5, 5, 2, -3, -4, 2, -20, 4, -10, 13, 15, -14, -7, -3, -8, 0, 5, 9, -8, -31, -9, 4),
    (6, 18, -3, -2, -27, 0, 12, -23, -12, -5, -34, 34, -32, 0, -2, -21, -14, 15, -40, -10, 4, -10, 22, 6, -42, -14, 23, -19, 22, 11, 26, 1, -2, -2, 20, -2, 14, 1, 7, -2, -15, 10, -11, 19, -23, 25, -8, -17, -12, 16, -34, -21, -4, -27, 6, -1, -29, 18, -30, 19, 29, 14, 9, -6, 16, -18, -4, 4, -12, -3, 25, 10, 9, 5, -2, 16, -15, -4, -17, 13, -3, 18, -23, 4, -5, 2, -4, -10, 12, -10, 18, -3, 5, 10, 21, -7, -5, -4, 0, -2, -2, 6, -3, -2, 7, -19, -8, 10, -2, 2, 2, -10, -12, 8, -6, -4, -17, 2, 11, -6, -2, -6, 7, 9, -3, -2, 26, 4, 1),
    (-7, 11, 14, 30, -30, 3, -10, -10, -37, -14, -48, -1, 29, 14, 23, -19, 7, 6, 8, -21, -28, 24, -19, -16, -34, -18, 1, 6, 6, 27, 1, 16, 4, -5, 13, -24, -4, -13, 12, -19, -20, -9, -13, -16, -6, 3, 13, -19, -34, 1, -6, -11, 19, -20, -16, -13, -31, -12, -18, -17, 17, 15, -11, -1, -6, 10, 2, 19, -25, 26, -18, -16, -45, -11, 30, 8, 1, 7, -14, -11, 6, 14, 12, -1, -22, -25, 18, -7, 4, 13, -6, -5, 10, 5, -3, 18, 0, -5, -3, -9, -14, 18, -17, 5, -9, 8, 3, 0, 18, 1, 5, -9, -8, 11, -8, -13, -8, -11, 2, -7, 1, -1, 6, -2, 10, -5, 11, 6, -25),
    (-49, -68, -10, -35, 21, -5, 16, 20, 23, 17, 34, 1, -12, 8, -17, 17, 7, -43, -20, 1, -14, -2, 14, 5, 20, 40, -26, -3, -15, -39, -7, -26, -24, 2, -24, -1, 0, 2, 10, -2, 15, -2, 0, 14, 13, -20, -6, 6, 23, 18, 1, -7, -25, 14, -15, 0, 5, 21, -3, 8, -19, -4, -8, -22, -10, 5, 5, 14, 25, -25, -7, 11, 22, 4, -14, -17, 10, -6, 4, 4, -4, -34, 7, -12, 2, 18, 9, -23, -6, 25, -13, -30, -28, -22, -7, -9, 14, -7, -1, -8, 20, -11, 0, 7, 17, 4, 3, -17, -13, -3, -4, 13, 11, -15, 1, 0, 20, 9, -14, 11, -2, 11, 0, -2, 0, 3, 9, -19, 2),
    (14, 16, -19, -7, 9, 7, -6, -24, -2, -27, 13, -14, 2, 18, -10, -7, -30, 15, 5, 18, 14, -13, -15, 31, 6, -1, 18, -18, 11, 5, 14, 22, 6, -14, 5, -11, -10, -8, -8, -7, -16, -18, 3, 9, 8, -1, -5, 2, -10, 4, 2, 7, 21, -3, 1, 5, -16, 2, 6, 11, 9, -5, 9, 11, 16, -6, 11, -14, -15, -4, 1, -20, -12, 2, -5, -2, -13, 10, 2, -4, -7, 16, -25, 6, -8, -5, -15, 11, -17, -8, 3, -7, 9, 9, -7, 11, 7, 11, -15, 6, -4, -6, -11, -8, 15, 3, 2, -4, -7, 14, 6, -8, -7, 2, -4, 2, 2, -6, 1, 5, -1, -2, 2, 4, 2, 7, 1, 10, -1),
    (-2, -40, 12, -46, -5, 14, -12, -38, 34, -19, 25, -1, -39, 11, 6, -17, 18, 8, -18, -10, 16, 5, 5, -21, 4, 11, -19, -4, 1, 19, 5, 14, 2, -13, -2, 1, -10, 2, -3, -12, 12, -5, 12, 14, 14, 6, 17, -18, 13, -16, -3, 0, -7, 16, 0, -4, -11, 15, 5, 12, -3, -28, 15, 7, -15, 10, -11, 22, 28, -14, 1, 14, 12, -14, -16, -12, 0, -12, 10, 16, 15, -17, 26, -29, 17, 25, -5, 1, -5, -1, -3, -39, -35, -3, -18, -6, 2, -2, -13, -7, 5, -8, -5, -2, 11, -5, -4, -11, -11, 0, 1, 9, 14, -16, 14, -19, 11, 22, -14, 3, -9, 14, -5, 1, -20, 7, -3, -10, 8),
    (-17, 6, 9, 0, 14, -31, 17, -9, -30, -22, 26, 26, -5, 6, 20, -26, 10, -6, 22, 12, -48, -2, 2, -25, 18, 26, -22, -2, -2, -4, -50, 33, -15, 17, -20, -4, -11, 4, 1, -6, -13, 19, 4, 16, -24, -19, 0, -17, 2, -6, 10, -32, -23, 7, -13, -18, 19, 18, 13, -16, -14, -23, -4, 8, -26, 4, 12, -7, -31, -6, -6, 17, -15, 14, 29, 17, -22, 5, -1, -7, -3, -2, -19, 13, -43, -30, -11, -14, 20, -2, 7, 7, 2, 17, 0, 30, -10, 3, 20, 17, 13, 6, 11, 35, -9, 0, -5, 8, -2, -21, 19, -2, -13, -5, 14, -2, -20, -12, -3, -3, 9, -2, -10, 7, -9, 5, 9, 9, 10)
  );
  ----------------
END PACKAGE CNN_Data_Package;
