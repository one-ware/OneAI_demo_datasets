library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.numeric_std.all;
use work.CNN_Config_Package.all;

PACKAGE CNN_Data_Package is
  CONSTANT Layer_1_Columns    : NATURAL := 128;
  CONSTANT Layer_1_Rows       : NATURAL := 128;
  CONSTANT Layer_1_Strides    : NATURAL := 1;
  CONSTANT Layer_1_Activation : Activation_T := relu;
  CONSTANT Layer_1_Padding    : Padding_T := same;
  CONSTANT Layer_1_Values     : NATURAL := 1;
  CONSTANT Layer_1_Filter_X   : NATURAL := 3;
  CONSTANT Layer_1_Filter_Y   : NATURAL := 3;
  CONSTANT Layer_1_Filters    : NATURAL := 12;
  CONSTANT Layer_1_Inputs     : NATURAL := 10;
  CONSTANT Layer_1_Out_Offset : INTEGER := 3;
  CONSTANT Layer_1_Offset     : INTEGER := 1;
  CONSTANT Layer_1 : CNN_Weights_T(0 to Layer_1_Filters-1, 0 to Layer_1_Inputs-1) :=
  (
    (24, -11, -25, -25, 8, -31, 30, 45, 64, 0),
    (18, 13, 64, -34, 20, 10, 10, 41, 33, -1),
    (-20, 27, -48, 40, 21, -53, 9, 32, -36, 0),
    (-23, 59, 49, -18, -7, 42, 17, 27, -32, -2),
    (-13, 24, -26, -31, 23, 49, -23, 0, -47, 1),
    (-51, -45, -5, 6, -9, 25, 48, 43, -16, -1),
    (44, 7, -4, 56, -20, -43, -29, -25, -36, 3),
    (22, -2, -4, 35, 13, 41, -16, -33, 53, 2),
    (19, -29, -62, 1, -15, -30, 34, 17, 18, -1),
    (24, -16, 1, 34, -19, -6, 25, 38, 7, -1),
    (-11, 36, 26, -46, -44, 28, -76, -39, 39, 0),
    (-17, 17, -15, 53, 43, -17, 2, 56, -1, -3)
  );
  ----------------
  CONSTANT Pooling_1_Columns      : NATURAL := 128;
  CONSTANT Pooling_1_Rows         : NATURAL := 128;
  CONSTANT Pooling_1_Values       : NATURAL := 12;
  CONSTANT Pooling_1_Filter_X     : NATURAL := 2;
  CONSTANT Pooling_1_Filter_Y     : NATURAL := 2;
  CONSTANT Pooling_1_Strides      : NATURAL := 2;
  CONSTANT Pooling_1_Padding      : Padding_T := valid;
  ----------------
  CONSTANT Layer_2_Columns    : NATURAL := 64;
  CONSTANT Layer_2_Rows       : NATURAL := 64;
  CONSTANT Layer_2_Strides    : NATURAL := 2;
  CONSTANT Layer_2_Activation : Activation_T := relu;
  CONSTANT Layer_2_Padding    : Padding_T := same;
  CONSTANT Layer_2_Values     : NATURAL := 12;
  CONSTANT Layer_2_Filter_X   : NATURAL := 3;
  CONSTANT Layer_2_Filter_Y   : NATURAL := 3;
  CONSTANT Layer_2_Filters    : NATURAL := 16;
  CONSTANT Layer_2_Inputs     : NATURAL := 109;
  CONSTANT Layer_2_Out_Offset : INTEGER := 3;
  CONSTANT Layer_2_Offset     : INTEGER := 0;
  CONSTANT Layer_2 : CNN_Weights_T(0 to Layer_2_Filters-1, 0 to Layer_2_Inputs-1) :=
  (
    (-12, 14, -5, 13, -27, -11, 28, 29, 1, 8, -21, 12, 23, 26, 20, -18, -7, -13, 23, -13, 18, -13, 4, -3, -9, -11, 15, -35, -6, 6, 20, -36, 10, 3, -21, 15, 0, 23, 12, -4, -26, -2, 4, 6, 16, 1, -3, 13, 5, -5, 36, 5, -11, -5, 20, -8, 19, -6, 8, 4, -2, -24, 15, -22, -2, -3, -8, -21, 26, 1, 0, 14, 17, 13, 27, 4, -19, 7, -9, 16, 3, 38, -15, 28, -19, 18, 16, 5, -12, -2, -2, -3, 6, 34, 17, 45, 14, -8, -11, -4, -10, -2, -18, -6, -20, -1, -5, 13, -4),
    (0, -26, -29, -1, 46, 12, -73, -29, -22, -11, 0, -27, -4, 0, -12, 11, 39, -10, -63, 7, -45, 27, 6, 14, 19, 33, -7, 28, 32, -19, -2, 17, -5, -3, 3, -4, 1, 14, -5, -11, 51, -8, -51, -11, -54, 13, -20, -14, 7, -13, -4, -13, 31, 8, -36, 13, -41, 1, -36, 20, 7, -6, 2, 1, 25, -8, -2, -3, -15, 20, -4, -5, 10, -18, -7, 12, 4, -9, -51, 6, -61, 10, -8, 11, 33, 33, 26, 18, 0, -5, -30, -17, -4, -2, -21, -5, 31, 23, -5, 20, 7, -4, -7, 27, -29, 31, -18, -13, 3),
    (-4, -5, 6, -22, -47, 17, -33, 6, 48, -8, -14, 17, 14, -1, 38, -10, -84, 29, -44, -36, 41, 23, -3, -26, 11, -14, 20, -31, -40, 35, -19, -34, 22, -35, 5, -21, 17, -27, -1, -26, 23, 5, -22, 8, 40, 1, -15, 22, -2, -23, 10, -33, -5, 23, -47, 4, 47, 38, -35, 38, 9, 25, 16, -23, -19, 27, -14, -20, 14, 13, -32, 14, 7, -15, 8, 19, 0, -30, -6, 26, 2, 15, 13, -5, 17, 25, -14, -14, 13, -9, -30, 15, -9, 16, 12, 20, -2, 19, -29, 5, -5, 11, -25, 29, 8, 13, 16, 16, -3),
    (-20, 4, 44, 27, -18, -15, 55, -22, 14, 14, -2, -17, 24, 25, -11, 20, -12, -41, 3, 2, -14, 11, 15, 33, 0, 18, -15, 15, 1, -33, -9, 19, -20, -3, 16, 27, 8, 10, 11, -2, 9, -18, 33, 6, -13, 2, -17, 3, -9, 37, 2, 8, -9, -19, 6, 23, -41, 16, -15, 12, 2, -13, -5, 26, -17, -9, -17, 13, -23, -3, -4, -8, -14, -6, 3, -2, -16, 2, 3, 26, 1, 16, 12, 28, -22, 14, 2, -5, -12, -7, 2, 9, -21, -16, -9, -1, -25, 10, 13, 12, -50, -17, -4, -15, -26, -14, 7, -9, -8),
    (0, -10, -5, -21, -26, 10, 22, 8, -18, 5, 13, 23, 7, -17, 19, 9, -26, 7, 25, -12, 29, -6, 2, 21, 7, 23, 19, 24, -9, -6, -4, 12, 25, -26, 7, 0, -18, -5, 3, 5, -34, 20, 20, 5, 25, -5, 0, 26, -32, 1, 11, -13, -33, 20, 19, -14, 40, 1, 38, 43, -12, -5, 14, 14, 15, 19, 31, 20, 35, -15, 23, 10, 28, 26, 14, -10, -8, 22, 6, -13, 18, -10, -12, -3, -8, 2, 24, 4, 6, 15, 3, 5, 39, -7, 34, 36, 12, -13, 10, 26, 31, 4, -14, -3, 41, 18, 40, 27, -5),
    (3, 31, -13, 21, 4, -43, -6, -1, -46, -24, 20, -3, -19, 29, 10, 18, 34, -45, -60, 28, 22, 3, 19, 14, 21, -13, 35, 2, 19, -3, -45, 0, 41, 20, -14, 1, -18, 7, -37, 22, 8, -17, -20, -25, -13, -1, 6, 0, -23, 0, -19, 13, 14, -21, -47, -3, -35, 3, 11, -14, 4, 3, 30, 15, 10, -11, -54, -5, 13, 4, -3, -20, -11, 18, -9, -24, 5, 62, 20, -13, 22, -21, 10, -36, -30, 0, -37, 9, -4, 2, -5, -7, -19, -30, 19, -27, -6, 14, -9, 24, -4, -17, -29, 26, -32, -13, -1, -23, -1),
    (9, -18, 5, -12, 22, -2, 12, 15, -1, -13, 18, -9, -16, 12, -27, -17, 1, -3, -13, -13, -42, -13, 32, -24, 16, -5, 4, 32, 19, -7, -34, 32, -47, -19, 36, 26, -28, 15, 15, -27, 21, 8, 14, -22, 2, -12, 11, 21, -20, 7, -22, 23, 8, -21, -31, -5, -39, 6, 8, -17, -10, 14, 10, 28, 8, 2, -37, 17, 15, 29, 27, 10, -24, 3, 18, -17, 23, -4, 22, -10, 12, -18, 18, -26, -7, -10, -12, -22, 11, -21, -54, 18, -9, -14, 38, 14, -13, 14, -10, 5, 0, -4, -29, 31, 0, 16, 22, 7, 0),
    (26, -17, -5, 18, 18, -47, 42, 8, 33, 9, 45, -26, -20, -6, -53, -29, -3, 5, 35, 15, -7, -38, -17, -45, 6, -14, -45, -19, -15, 24, 6, 11, 31, -14, -3, -36, -1, -1, -30, -4, -42, 7, -6, 14, -4, -27, -23, -32, 16, -17, -42, 6, -21, 28, -14, -22, 5, -18, -12, -20, 40, 5, -38, 14, 14, 28, -38, 11, 36, 21, 4, 24, 3, 14, -6, 26, -7, 12, -20, -15, -10, 5, -12, 23, 26, -7, -22, 25, -6, 25, -15, -7, 7, 9, 4, 3, 31, 12, -32, 5, 14, 37, 5, 35, 9, 12, -9, -7, 0),
    (19, -7, 23, -6, 19, -9, 17, 14, -6, 9, 8, 35, -9, -3, 13, 37, 3, -32, 47, -12, -21, 23, 0, 7, -2, 21, -2, 19, -3, 4, 43, -18, -31, 12, -28, 16, -35, -10, 2, -9, 46, -17, 23, 0, 18, 1, 15, -28, -4, -18, -49, 1, 7, 20, -1, 15, 22, -40, -23, -15, -2, 4, -12, -32, -16, 20, 14, -32, 19, -29, -21, -36, 12, 16, -36, -41, -17, 27, -43, 18, -15, 3, -24, -24, 5, 1, -6, -21, -21, 15, -52, -14, 14, 10, -23, -1, 20, -1, 1, 17, -8, 9, -57, 28, 35, 5, 0, 30, 0),
    (6, 33, 7, -10, -18, -14, 21, 23, 3, 36, -18, 15, -4, 4, -11, 22, -39, -10, 23, 9, -21, 16, -7, 19, 15, -5, 0, 9, 15, 14, 12, -2, 10, -7, -12, -10, -1, -7, 2, 17, -24, 15, 29, 20, 0, 28, -10, 15, 4, 10, -15, 15, -21, 0, 7, 13, 0, -12, 9, 27, -4, 9, -20, 16, -3, 8, 24, 15, -13, 2, 13, 2, -4, -20, -6, 26, -17, 22, 28, -1, 20, -2, -8, 1, 14, -11, -26, 15, -19, 16, 25, 7, -1, -17, -28, 11, 4, 6, -12, 15, 9, -15, 10, -5, -13, 1, 17, 26, -3),
    (11, -7, 26, -22, 36, 31, -13, 47, 38, 29, 10, -5, 20, -43, -25, -14, -55, -6, -17, -8, -8, 17, 12, -13, 2, -10, -53, -4, 8, 19, -8, 27, -46, 14, 10, -27, 23, 3, 40, -11, 8, 48, 21, -12, 41, 38, 20, -10, -23, -38, -3, -48, -127, 16, 15, -25, 1, -18, -21, 11, 2, 0, -43, -18, 11, 9, -33, 16, -28, -21, 28, -12, -3, -19, -2, 6, -34, 24, 28, 2, 33, 16, -33, 13, -19, 1, -5, -28, -69, -36, 37, 10, -14, -31, 3, 1, 22, 22, 11, -18, 17, -25, -18, -2, 18, -15, 1, 2, 6),
    (1, -6, -18, -9, -11, 21, -3, 4, -14, -32, 6, -5, -37, 8, -25, 24, 1, -16, -6, -19, 9, -30, 54, -27, -31, 24, -11, 40, 5, -47, 13, -24, -22, -19, 36, -29, 23, -19, 9, -24, -57, 46, -26, 12, 24, 16, -26, 27, -3, -11, -1, -23, -61, 24, -32, -11, 42, -17, -31, 17, -6, -26, 4, 0, -9, -5, -19, -25, 17, 4, 22, 3, 13, 2, 25, -5, 31, 17, -7, 9, 16, 35, -1, 30, 0, -3, 46, -5, 18, 19, -39, 13, 43, 30, 9, 7, -5, 0, 23, -16, 15, -14, -20, 1, 18, 14, 9, 12, 0),
    (-21, -40, -14, 6, -19, 8, -4, -34, 36, -4, 5, -13, 18, 21, 6, 1, -30, -16, 11, 11, -32, -34, 8, -7, 2, -3, 17, 19, -7, 5, 23, -13, 13, -7, 16, 10, 16, 8, 17, -13, 2, -22, 21, 13, -4, -15, -13, -18, 13, 3, 14, -21, 2, -33, -25, 24, -6, -11, 25, -16, -9, -19, 19, -17, 11, -25, 25, -5, 32, -2, -42, -25, 22, -23, -9, -37, -5, 23, 26, 11, -2, 32, -6, -25, -25, 21, -24, 23, 37, -11, -14, -11, 33, 16, 20, -16, -16, -36, -14, -17, -11, -22, 41, -38, 3, 14, -31, 8, 4),
    (10, -20, -5, 18, 18, 18, -30, -6, -15, 27, 4, 8, 33, 0, -4, 14, 33, 7, -13, -12, -4, 4, -16, 11, 27, -15, 22, -8, 28, -12, -26, -24, -3, 20, -33, 11, 8, -12, 25, -1, -1, -21, -38, -13, -31, 22, -27, -12, 30, 21, 26, -17, 26, -25, -34, -2, -4, 0, -33, 9, 19, -12, 9, -2, 13, -29, -28, -8, -25, 7, -33, -4, 37, 22, 28, 9, -32, -23, -23, 8, 7, 28, -14, 23, -1, 33, 26, -12, 1, -26, -19, 10, 16, 36, -7, 26, 6, 1, 32, -23, 3, -18, -38, -27, 10, 35, -19, -4, 4),
    (19, 40, 11, 25, -7, 3, 35, 26, -37, 22, 26, -11, 2, -3, 45, 38, -9, -25, 27, 19, 13, 16, 32, 22, -27, 22, 28, -14, -17, -52, -2, -12, 36, -10, 14, 20, 14, 2, 22, 15, -5, 18, 56, 2, 1, -11, -16, 9, 1, -6, 20, -1, -24, -16, 31, -25, -18, 19, -27, 11, -30, -24, 12, -20, -35, -36, 13, -24, -4, 8, 5, 12, -18, -28, 21, -18, 24, 12, 26, -3, -6, -11, -7, 5, 7, -24, -5, -17, -23, -12, 15, -20, -18, -22, -20, -27, -4, -20, -53, 18, 0, -25, 3, -19, -25, -5, 10, 10, -4),
    (-16, 15, 15, 12, 37, -22, -13, 8, 24, 1, 7, -7, 22, 19, -6, 6, 37, -9, 2, -4, 11, -16, 35, 22, 36, 12, -3, 36, 14, -3, 9, 40, -16, 25, 9, -7, -29, -7, -14, -9, 50, 0, -17, -34, 38, -32, 2, -35, -34, -1, -40, -18, 20, -21, -14, -11, -18, -16, -3, -21, -6, 0, -43, 20, 9, 12, 29, 4, -10, -19, 4, 14, 3, 18, 25, 18, -82, 28, -40, -15, 22, 29, -21, 0, 0, 11, 10, -31, -59, 33, -59, -35, 27, -13, -42, -4, 2, -20, -24, -15, -11, 39, -33, -22, 37, -6, -20, -4, 1)
  );
  ----------------
  CONSTANT Layer_3_Columns    : NATURAL := 32;
  CONSTANT Layer_3_Rows       : NATURAL := 32;
  CONSTANT Layer_3_Strides    : NATURAL := 2;
  CONSTANT Layer_3_Activation : Activation_T := relu;
  CONSTANT Layer_3_Padding    : Padding_T := same;
  CONSTANT Layer_3_Values     : NATURAL := 16;
  CONSTANT Layer_3_Filter_X   : NATURAL := 3;
  CONSTANT Layer_3_Filter_Y   : NATURAL := 3;
  CONSTANT Layer_3_Filters    : NATURAL := 24;
  CONSTANT Layer_3_Inputs     : NATURAL := 145;
  CONSTANT Layer_3_Out_Offset : INTEGER := 3;
  CONSTANT Layer_3_Offset     : INTEGER := -1;
  CONSTANT Layer_3 : CNN_Weights_T(0 to Layer_3_Filters-1, 0 to Layer_3_Inputs-1) :=
  (
    (-36, 55, -38, 15, -3, -72, -14, 113, 33, -31, -28, -30, -23, 28, 60, -31, -1, 38, -15, 37, -18, -55, 6, 64, 48, -37, -4, -34, -53, 17, 67, -77, -27, -16, -11, -18, -10, 18, -26, 24, 19, 30, -36, 22, -42, 25, 15, 3, 19, 71, 10, 31, 47, -62, -14, 102, 75, -28, -38, -11, -37, -10, 90, -25, 27, 51, 20, 32, 36, -47, -12, 95, 38, 30, -29, -1, 20, 11, 63, 0, -25, -38, -10, 11, -46, -4, -60, 9, 35, -17, -8, 3, -19, -3, 19, -13, 12, 14, 24, 41, 39, 6, -5, 52, 61, -34, 35, -13, -40, -39, 20, -32, -51, -32, -6, 24, -53, -31, -55, 50, 58, -31, -3, 23, -49, -72, 3, 50, -33, -56, 24, -35, -94, -31, -105, -18, -11, -34, -40, 56, -12, -31, -1, 91, -4),
    (-66, -18, 9, -63, -1, -37, -4, 52, 51, 7, -26, -38, -12, -62, -52, -18, -12, -69, 14, -31, 30, 39, -36, -13, -7, -59, -7, 48, 7, 18, -36, 36, -55, -37, 27, -57, 37, 75, -5, -44, -7, 1, 17, 71, 3, 9, -53, 37, -48, -20, -79, -32, -1, 4, 10, 15, -25, -38, 89, -28, 30, -24, -24, 11, 8, 11, 19, 28, 10, 17, 28, -50, -12, -42, 82, 92, 14, 13, 18, 58, -6, -33, 43, -16, 25, 36, -5, -68, -14, 4, 26, 80, -4, -3, -19, 60, 19, -16, -44, 1, -38, 55, 42, -3, -20, -40, 47, -8, -22, -18, -60, -15, 41, 46, -1, 14, 8, 2, 85, -19, -39, 43, 109, 41, -34, 61, 4, 7, -3, 31, 26, -16, -8, -11, 18, -36, -42, -35, 45, 37, -44, -23, -16, 20, -3),
    (-3, -17, -23, -29, -29, -53, 17, 16, 9, -30, 15, 34, -11, 15, 15, 10, -44, 4, 46, 16, 0, -88, -34, 38, 4, -6, 25, 30, -21, 29, -4, 21, -3, -14, 62, 17, -18, -48, -6, 44, 24, 76, -34, 15, -83, 39, -28, 15, -39, 35, -18, 21, 1, -28, 42, -21, -13, 20, 21, -18, 18, 21, -26, -55, -31, -3, 50, 11, -6, -51, 7, 43, 80, -43, -46, 2, -34, 34, 44, -32, -10, 48, 51, 2, -47, -41, 3, 57, 77, 39, -54, -15, -35, 36, 14, -4, -30, -54, -93, -9, -2, 8, 3, -41, 36, -51, 28, -9, -2, -67, -69, 25, -52, -58, -71, 40, 8, -32, -37, 34, 91, -23, -49, -13, -5, -44, 25, -10, -52, -52, -18, 43, -2, -15, -41, 37, 56, 50, -56, 2, 10, -52, 22, 39, 2),
    (46, -24, 55, 19, 18, -46, -46, 37, 57, 19, 32, -11, -36, -12, 69, 47, 42, 36, 4, 45, 53, 11, -7, 40, 63, 45, -29, 20, -10, -19, 31, 22, 35, -44, -48, 15, -44, -48, -16, -66, 41, -14, -7, 3, -26, -47, -11, 2, 1, 7, 25, -41, -5, -24, -73, -5, 43, 3, 28, 11, 48, -5, 20, 57, 16, -42, 12, -40, -45, -1, -103, 48, 54, -51, 0, 23, -17, 3, 16, 48, -1, -72, -28, 6, -52, -29, -78, 28, 44, -65, -23, 52, -15, 22, 24, -36, -10, -32, 39, -48, 14, -44, -100, 26, 87, -48, 3, 65, 49, 1, -8, 27, -38, 6, 46, 18, 14, -96, -52, 73, 57, -20, 24, -9, -32, 37, -11, -48, -53, 32, 25, 20, 33, -25, -44, 9, 57, -23, 64, -8, 36, -4, -57, -22, 10),
    (-17, 24, 7, 17, -30, -4, -42, 15, -7, -3, -22, -10, 23, 33, -16, -54, -21, -29, 63, -17, 8, -44, -65, 25, 4, -7, -59, -15, -15, 6, -5, -47, -46, -91, 39, -9, -39, -54, -51, 37, 65, 41, -33, 14, -39, -47, 0, 31, 33, -20, 22, 7, -3, -51, -24, -7, -39, -1, 48, -12, -4, 51, -43, -48, 23, 12, -26, -42, 9, -32, -21, -13, 3, 17, 3, -26, 66, 27, -45, -89, -14, -34, -5, -11, 35, -65, 2, 13, 25, -34, -26, -13, 25, 31, 17, -37, 39, 37, 24, 56, 21, -12, 21, -22, -23, 3, 7, 6, -14, 42, 23, -6, 47, 35, 1, 0, 7, -16, -10, -32, -29, 16, -19, -15, 24, 35, -21, 15, 9, 55, 26, 46, 6, -17, -5, 55, 25, -12, -18, -14, 7, 65, 7, -27, 4),
    (-4, 10, 7, 3, 37, 19, -55, 6, -22, 5, -29, 8, 17, 66, 8, 34, 33, 43, 16, 8, -5, 46, -17, -11, 5, 38, -54, 35, 2, -25, -13, 57, 29, 32, 29, 23, 34, 9, -3, 4, 7, 21, 10, -11, -13, -15, -54, 36, 31, 1, 20, 24, -9, -7, -44, 10, -3, -28, -28, 51, -16, -31, -6, 17, 33, 28, 14, 36, -36, 38, -72, 19, 29, 50, -42, 20, -9, -12, -36, 80, 25, 21, 50, 49, -25, 30, -4, 9, -12, -20, -43, 52, -78, -1, -67, 11, 3, -5, 12, 34, -31, 23, -34, -27, 10, 8, -79, -6, 0, -70, -17, 25, -6, 3, 48, 52, -26, 77, -54, 26, 14, 21, -12, 39, -62, -63, -19, 35, 14, 19, 4, -4, -12, 47, 12, 24, -5, 31, 30, -6, -51, -40, -53, 14, -4),
    (14, 4, 15, 15, -4, -12, 0, -27, 5, 45, -12, 64, -10, -2, -23, 5, 45, -3, 34, 14, 46, 23, 23, -37, 12, -31, -12, 60, -66, -9, -15, 28, -34, -8, 8, 37, 21, 43, 38, -21, 7, 2, -2, 48, 10, 34, 7, 33, -1, -45, 44, 15, 14, 21, -19, -33, 4, 0, -7, 76, -19, -20, -34, 45, -8, -68, 81, 12, -4, 66, -30, -34, 0, 52, -70, 117, -56, -21, -62, 75, 34, 5, 19, -25, 22, 70, -4, -39, 7, 34, -37, 53, -45, -28, -47, 83, -28, -5, 40, -32, 18, 58, -9, -54, -3, 44, -11, 82, 20, -28, -24, 70, -7, -26, 40, 7, 47, 59, -28, -3, 9, -13, -26, 60, -13, -38, -55, 50, -28, -34, 36, 36, -1, 28, -50, 7, 2, -44, -27, 36, -4, -38, -27, 12, -5),
    (36, 64, -29, 37, -3, -56, 10, 41, 24, -8, -7, -34, -35, -10, 62, -11, -4, 90, -41, 10, 18, -46, 44, 9, -40, -13, -3, -58, -2, 13, 61, -31, 12, 57, -41, 68, 16, -13, 64, -18, -46, 9, 22, -25, 21, -8, 6, 2, -2, 35, -44, 19, 28, -58, 41, -18, -3, -6, 42, -88, 12, 14, 56, -2, -29, 60, -76, -8, 2, -49, 65, -5, 14, -15, 59, -58, -7, 52, 63, -37, -7, 26, -83, -6, -16, -36, 30, -36, -20, 14, 27, 5, -17, 17, -1, 17, -18, 16, -59, 20, -2, -31, 47, -14, -5, 6, 39, -39, -47, 18, 0, 9, 46, 22, -87, -9, 3, -23, 54, -26, 19, -44, 68, -17, 52, -2, 4, 18, 14, -14, -37, -16, -23, -42, 32, -71, -38, -27, 5, 57, 27, -10, 18, 15, -2),
    (3, -11, -40, -1, -37, 20, 41, -48, -88, -71, -38, -33, 16, -75, -102, -25, 31, 29, 14, 14, -39, 20, 26, 8, 1, 4, -39, -43, -36, -38, 9, 4, 15, 54, -3, 26, 17, -33, 9, 60, 83, 71, -9, -44, -75, -8, -2, -15, -29, -20, -59, -1, 1, 37, 34, -12, 53, -18, -54, 53, 10, 17, -70, 73, -51, -60, -53, -7, -47, -40, -29, 8, 86, 28, -31, 44, -29, 18, -61, 72, -50, -73, -1, 17, 24, -51, -9, 51, 54, -23, -51, 1, -68, -5, -23, -13, 5, -20, 29, -35, 5, -43, -29, 16, -4, -7, 4, 61, 99, 0, -66, 22, 20, 9, 51, 8, 39, -37, -32, 2, -17, -13, -67, 29, 13, -15, -19, 81, 26, 23, 65, -46, -25, 39, -20, 37, 59, -40, -26, 39, 31, 25, -36, -2, 1),
    (-27, -9, -14, -21, 34, -65, 34, 2, -28, -20, 68, -55, 12, -6, -47, -4, -5, 46, 11, 46, 46, 31, -3, -7, 24, 10, 93, 6, 42, -23, 38, 53, -48, -27, -25, -44, -39, 64, -27, -80, 12, -61, -6, -36, -45, -14, 2, -62, -35, 19, -18, 11, 46, -36, 56, 7, 13, -49, -23, -33, 8, 0, -96, 22, 48, 31, 38, -5, 23, 14, 32, -28, 7, 24, 54, 3, -9, -35, 55, 49, -57, -32, -45, 15, -82, -43, -66, -36, -36, 13, 5, 7, 4, -40, -25, 22, -24, 17, 12, -46, -18, 1, -44, -24, -52, -36, -36, 35, 42, -23, -86, 60, 28, 23, 5, -27, 33, 3, 75, 17, -1, 3, 81, -24, -7, -56, 25, -7, -10, -60, -26, 28, 6, -54, -8, -23, -66, -41, 32, -20, -33, -4, -12, 20, 0),
    (26, -12, -31, 37, -2, -13, 0, 23, -11, -30, -16, -33, -36, -46, 17, -6, 39, -2, -54, -20, -9, 15, -24, -9, -13, 14, 25, -65, -10, -48, 22, -46, 11, -18, -32, 16, 50, 1, 1, -5, 20, -32, -30, -34, 16, -21, -17, -16, 31, 5, -63, 25, 56, 18, -6, -8, -16, 12, 1, -54, 11, -37, 23, -12, 34, 6, -54, -9, 87, 54, 7, -42, -68, 41, -2, -83, 47, -18, 5, -11, 63, -7, -30, 45, 28, 30, 7, -8, -6, -14, 12, -46, 31, -17, -39, -15, -8, -22, -1, 13, 28, 5, -50, 30, 13, 25, 18, -18, -31, -23, 10, -11, 59, -13, -11, 57, 46, 11, -4, -18, -1, 0, 7, -52, -14, 7, -17, -20, 11, 28, -17, -10, 75, 12, 12, -29, 32, 34, -10, -11, -48, 22, -53, 7, -14),
    (46, 0, -17, 2, -25, 1, 24, -2, 8, -18, 15, -38, -69, 27, 59, -1, 12, 60, -3, 61, -34, -31, -10, 40, 64, 65, -27, 0, -96, -1, 82, -1, -22, 28, 1, 71, 30, -28, -31, 50, 72, -8, -2, 5, -31, 2, 64, 9, -59, 26, -4, 33, -39, 32, -19, -4, 41, -34, -25, 67, -3, -17, -2, 48, -66, -21, 17, 8, -35, -19, -30, 55, 80, 56, -96, 39, -27, -55, 1, 27, -18, -40, -35, 65, 35, -32, -32, 92, 88, 35, -67, -41, -13, 7, 12, 6, -23, 2, 1, 4, -62, -59, -40, 29, 5, -46, -36, 16, 28, -33, -42, 80, -13, -25, 39, -50, -75, -62, -46, 35, 30, 31, -62, 20, -10, -15, -29, 27, 0, 0, -5, -49, -22, -27, -15, 26, 7, -8, -60, -27, -41, -7, 22, -73, -8),
    (33, 57, -63, -28, -28, -38, 43, -15, -33, 30, -5, -39, 24, 2, -16, -2, -1, 26, 18, 21, -16, -23, 11, -2, -11, 29, 24, -4, 3, -26, -35, 17, 25, 57, 22, 57, 24, -8, -52, 52, 32, 25, -89, -22, -72, -33, -29, -7, 38, 48, -52, -34, -45, 21, 52, -84, -30, 23, 36, 66, 39, -21, -63, 36, 56, 20, 40, 10, 58, 66, 5, -63, -11, 9, -11, 73, -55, 20, -107, 37, -43, -8, 75, 16, 48, 16, -50, 20, 20, -2, -65, 27, -99, -17, -64, 28, 2, 30, -8, -44, -24, 25, 13, -41, 5, -20, 17, 87, -1, -47, -43, 42, -36, -4, 30, -33, 17, 102, 7, -36, -39, -22, 5, 99, 9, -11, -91, 44, -13, -57, 22, 37, -14, 26, 32, 20, 9, -42, -10, 50, -4, -23, -56, 26, -4),
    (-37, 6, 3, 24, 37, -46, 55, 27, 21, 39, 60, -36, -13, -6, 67, -14, -7, -17, -93, 48, 0, -60, -67, 12, 16, 1, 20, -59, -41, 41, 1, -53, -50, -29, -55, -57, -87, -90, -109, -49, 15, -10, 19, -4, -39, -11, -36, -35, 6, 30, -103, 48, 0, -97, 44, 45, 15, 7, 38, -102, -3, 36, 59, -51, 41, 32, -70, 32, -51, -56, 32, 22, 7, -32, 48, -116, 15, 7, 8, -116, -10, 35, -7, -6, -9, 9, -15, 22, 19, -53, -16, -54, -25, -27, -35, -124, -28, -27, -77, 44, 0, -89, -18, -30, -42, 27, -18, -16, 6, 7, 36, -61, -2, 45, -45, 46, -28, -5, 66, 5, -47, -42, -7, 5, -5, 13, 14, -24, -11, -43, -47, -12, 30, 31, 56, -34, -37, 5, -54, 10, -2, 14, -7, 57, -4),
    (-84, 5, 7, -43, 9, 17, -27, -36, 31, -43, -59, 23, -22, -60, -37, 35, -26, -56, -51, -21, -1, 15, -4, 20, 73, -36, -14, 20, -31, -10, -76, 35, -32, -39, 15, 17, -11, -28, 13, 14, 34, 13, -78, 49, -14, 28, -43, 47, -49, 3, 21, -43, -2, -22, -38, 13, -5, 8, -51, 60, 30, 12, 21, 40, 29, -38, 60, -11, 24, -1, -26, 19, 38, -8, -44, 104, 30, 27, -38, 80, 4, -20, 52, 0, 38, 28, -40, 37, 62, 35, -31, 87, -42, 24, -58, 78, -1, -9, 7, -3, 32, -31, -5, 11, 28, -9, 26, 18, -18, -1, 8, -37, 0, -10, 47, -14, -16, -25, 0, -28, 2, -28, -4, 76, -24, 14, -30, 34, -32, 31, 35, 24, -2, -3, -23, 5, 14, 6, -28, 62, -22, 31, -53, 45, -2),
    (-6, -9, 23, 38, -21, 21, 19, -58, 11, 51, -37, 62, -23, 13, 25, 17, -11, 26, 2, 4, 32, 106, 27, -64, -27, 35, 20, 57, 33, 5, -23, 37, 33, -20, 16, 42, -5, 75, 18, -52, -68, -30, 37, 64, 64, 2, -39, 39, -10, 19, -45, -2, -29, 79, 20, -65, 6, -39, -31, 30, -11, -29, -3, 47, 1, 13, -21, 23, -37, 98, 33, -111, -49, -23, 23, 28, 69, 4, 11, 18, 2, 23, -10, 28, 0, 21, 29, -127, -54, 48, 55, 3, 37, -34, -13, 34, 15, -10, 25, 9, 3, -78, 16, 2, -39, 13, 32, -10, 29, -9, -37, 24, -29, 17, -38, 18, -32, -4, -2, -52, 25, -76, 10, -19, -10, -31, -70, 23, -69, -66, -25, 7, -75, 7, 19, -96, 34, -22, 19, 10, 43, -5, -37, -17, 3),
    (9, -69, 10, 18, 17, -18, 10, 11, 9, 1, 25, 1, 17, -45, 27, 32, -26, -88, 17, -26, 57, 27, 39, 3, -19, -20, -39, 4, -6, -17, 61, 14, 1, -38, 24, 27, 69, 31, -6, -14, 24, -37, -13, -20, -71, 1, 16, 18, 4, -37, 28, -7, 59, 22, -7, -7, -23, 8, 2, 47, 1, -22, 38, 2, 42, -86, 32, 20, 64, 29, -29, 8, 27, 3, -33, 38, -31, -49, 46, 2, 15, -45, 41, 26, 62, -5, -7, 5, 28, 49, -46, 46, -4, -42, 1, 27, 28, -34, 23, -14, 23, 6, -2, 7, -8, -44, 31, 12, -15, -6, 12, -17, 4, -39, 32, -9, 61, 7, -4, -8, 8, 36, 9, 16, -50, -28, 13, -3, 28, -15, 7, -9, 16, 7, -50, 4, 22, -17, -16, 24, -32, -26, -5, 17, -12),
    (33, 11, 1, -32, -33, 36, -36, -8, -36, 45, 32, 0, -13, 0, -79, 16, -46, -47, 42, -36, 1, 116, -3, -96, -45, -43, 7, 36, 61, -11, -54, 58, 1, -59, -1, -28, -60, 55, 23, -47, -7, -18, 30, 48, 71, -31, -84, 71, 41, 49, 42, 14, -20, 28, 64, -67, -68, 14, 49, 24, 65, 38, -26, -33, 32, 40, -14, -24, -13, 72, 40, -53, -71, 25, 57, 17, 55, 23, -52, 30, 15, -9, -24, -35, -37, 101, 54, -75, -71, -60, 18, 29, 8, 25, -22, 56, 14, 35, 11, 41, 28, 37, 88, -55, -46, -40, 65, 5, 20, 56, 14, -10, 14, 27, -3, 17, 48, 61, 115, -41, -82, -46, 67, 29, 47, 49, 10, 9, -25, -19, 23, 35, 39, 59, 28, -35, -25, -38, 24, 12, 63, 67, -2, 6, 7),
    (1, 11, 39, -23, 6, 11, -62, -1, 59, -35, 3, 19, -31, -71, -17, 0, -58, 6, -36, -47, 61, -38, 13, 29, 22, -31, -10, -48, 33, -34, -25, -13, 59, 2, -39, 69, 30, -29, 59, 27, 18, -15, 56, -16, 4, 28, 32, 12, 9, 28, -6, -70, -7, -9, 4, -31, -18, -49, -11, -14, -42, -14, -24, 40, -50, -36, -27, -49, -32, -41, 13, 5, 8, -18, 62, 46, -13, -25, -62, 26, 40, -6, -39, 54, 43, -7, 91, 2, 4, 35, 103, 53, 4, 44, 9, 51, 43, -55, 25, -15, -40, 41, 68, -72, 2, -39, 48, -11, -2, -7, -53, 55, 1, -16, 0, 28, -4, 26, 56, -14, -15, -39, 44, 35, 41, -55, -81, 56, -9, 52, 1, 13, 34, 29, 71, 3, -23, 25, 76, 54, -18, 31, -13, 35, -12),
    (-12, 33, 5, 27, -37, -45, -43, 0, 20, 9, -12, 2, -5, 34, -16, -9, 29, -28, 27, -7, 0, -17, 10, 2, 4, -14, -64, -16, -32, -28, 16, -18, -23, 30, 31, 4, -15, 20, -28, -12, -9, 3, -24, -16, -18, 26, 20, -23, 6, 4, -20, 63, -1, -52, -3, 25, -21, 21, -16, -24, -12, -8, 31, -69, -24, -24, -13, -5, -16, -26, -49, 31, -7, 48, -18, -21, -48, 43, 50, -26, -8, 38, -6, 35, 38, -20, -25, 15, 5, 14, -16, -33, -61, 30, 8, -39, 27, 50, 20, -4, 2, -24, -36, -21, -27, 12, 23, 1, 2, 47, 30, -30, 48, 17, -2, -1, 17, 18, -17, 9, 14, 31, 1, -28, -34, 2, 11, -21, 40, 51, -12, 16, -34, 3, -21, 31, -19, 23, -20, -3, 10, 18, 13, -24, -8),
    (-21, 70, -45, 0, -12, 51, 13, -38, 24, -16, -14, 25, 32, 17, 5, 29, -14, 61, -85, 8, 25, 75, 30, -113, -6, -24, -12, 77, 85, -32, -12, 62, -20, 54, 59, 47, 10, 57, 27, -56, -33, 33, 54, 96, 41, 4, -13, 48, -28, -4, -87, -40, -45, -81, 22, -6, 43, -49, -45, 11, 4, 11, 8, -44, -79, 34, -24, -23, -6, -24, -13, -29, 100, -30, 20, -9, 49, 9, -2, -10, 4, 2, -14, -11, -48, 14, 22, -5, 41, 1, 10, 47, -50, -41, -62, -11, -58, 5, 19, -18, -35, -36, -67, 59, -18, -19, -72, -10, -64, -14, -79, 11, -28, 24, -1, 12, -7, -52, -46, 55, 11, 5, -10, -22, -43, -4, -1, -81, -8, -8, 6, -32, -27, -87, -6, 10, -3, -10, -37, -36, -50, -17, 36, 8, 13),
    (29, -8, -17, -3, 15, -57, -4, 17, -32, 5, -24, -39, -22, -55, 18, -74, -9, -42, -32, -37, 23, 0, 33, -10, -40, 26, -17, 6, 14, 8, 9, -65, 10, -6, -22, 39, -4, -5, 56, 15, 14, 22, 2, 1, -18, -75, -27, -30, 18, -55, 41, 19, 39, -26, -2, -5, -35, 51, 30, 4, 25, -44, 0, 0, 29, -50, 50, 51, 29, 41, 11, -51, -27, 55, -23, 15, -10, -43, -43, -1, 39, -19, 10, 63, 35, 8, 32, -10, -27, 45, -56, 0, -43, -42, -29, -19, 40, -27, -27, -8, -12, -6, -17, 9, 9, 48, 27, -29, -60, -30, -7, -33, 28, -18, -7, 39, 36, 1, 2, -19, -44, 29, -32, -15, 13, -27, -40, -23, -22, 15, -7, 41, 36, -40, 66, 54, 24, 25, 6, -10, -27, 28, -70, 0, -6),
    (27, 7, -2, -21, 27, 22, 15, -34, -22, 19, 25, 4, 32, -33, -5, -27, -8, 5, -43, -24, 19, -1, -13, -54, -52, 21, 6, -6, -34, -27, 0, 21, 9, 22, -13, -25, 23, 36, -45, 8, 2, -27, -23, -1, -37, 30, 11, -29, -25, -15, -4, 23, 53, 9, -17, -11, 6, 62, 28, 16, -26, 20, 4, -11, 72, 17, -41, -22, 50, 12, -17, -45, -30, 93, -3, -28, 22, -91, -52, 1, 42, 24, -13, 4, 13, 26, 8, 10, 51, 30, -28, -47, 12, -21, -49, 4, 41, 16, -10, 60, 2, -27, -8, 53, -22, 21, -34, 0, -10, 2, -17, 18, 50, 18, 1, 30, 42, -24, -28, 4, 4, 46, -27, -13, 1, 40, -42, 13, 9, 13, 5, -17, -10, -16, -29, 31, -5, 53, -31, -12, -15, 1, -43, 20, -12),
    (0, -22, 13, 34, 1, 104, -63, -29, -54, 33, 91, -40, 33, 51, -10, -23, -40, -72, 8, -51, -38, -3, -44, 15, 52, -28, 24, -4, 16, -35, -47, 1, -69, -51, 53, 40, -46, -53, -26, 11, 43, 47, -54, -39, 16, -20, 4, 13, 44, 20, 20, 38, -4, 87, 15, -64, -42, 43, 77, -18, 93, 58, -5, -49, 28, -8, 8, -19, -2, 33, -40, -89, -40, 20, -21, -16, 27, -27, -24, -23, -76, -28, -31, -53, -60, -10, -70, -32, 27, 20, -41, -20, 12, -43, -3, 53, 72, 12, -27, 39, 56, 1, 87, -70, -28, -25, 64, -6, 52, 22, -31, -5, 43, -9, -28, 31, 22, 14, 13, -65, -80, -11, 9, -10, 0, 41, -24, -63, 9, -33, -7, -55, -32, 16, -50, -62, -20, -2, 19, 17, -20, -54, -12, -14, 4)
  );
  ----------------
  CONSTANT Layer_4_Columns    : NATURAL := 16;
  CONSTANT Layer_4_Rows       : NATURAL := 16;
  CONSTANT Layer_4_Strides    : NATURAL := 2;
  CONSTANT Layer_4_Activation : Activation_T := relu;
  CONSTANT Layer_4_Padding    : Padding_T := same;
  CONSTANT Layer_4_Values     : NATURAL := 24;
  CONSTANT Layer_4_Filter_X   : NATURAL := 3;
  CONSTANT Layer_4_Filter_Y   : NATURAL := 3;
  CONSTANT Layer_4_Filters    : NATURAL := 32;
  CONSTANT Layer_4_Inputs     : NATURAL := 217;
  CONSTANT Layer_4_Out_Offset : INTEGER := 3;
  CONSTANT Layer_4_Offset     : INTEGER := 0;
  CONSTANT Layer_4 : CNN_Weights_T(0 to Layer_4_Filters-1, 0 to Layer_4_Inputs-1) :=
  (
    (18, 6, 1, 3, 0, -6, -23, 25, -5, -7, 22, -15, -22, 22, -1, -23, -14, -9, 17, 16, -10, 0, 17, 27, 24, -3, 13, 24, 11, -14, -5, 27, -16, 2, 3, 5, -31, 10, -8, -20, -13, -12, 33, 1, -33, -14, -4, 7, 17, 4, 5, 32, -15, -2, -12, 11, 1, 20, 3, 19, -16, -2, 9, 13, 10, -4, 13, -21, 8, 5, -16, -9, 1, 12, 3, -13, 13, -6, 12, 19, -10, 19, 19, -13, 5, 3, -53, 6, -18, 5, 10, -12, 10, 13, -12, 16, -12, -7, -10, 4, -21, -11, -7, 23, -7, 10, 5, -11, 13, 8, -29, 19, -10, -15, 29, 0, -13, -6, 14, 16, 11, -14, -4, 19, -21, -15, 8, 4, -2, 25, -29, -2, -27, 1, 24, 2, -5, 6, -18, -22, 5, 6, -22, 1, -19, 7, -16, -20, -13, 25, 21, 1, -19, 1, 19, -13, 16, -15, -52, 16, -5, -6, 2, -24, 8, -14, 5, 17, -2, -13, -2, 5, -5, 5, 18, -8, -20, -3, -12, -16, 25, -23, -26, 16, -2, -23, -39, -1, 22, -10, 0, 17, 5, -15, 2, -20, -21, 8, -5, -18, -19, 15, -23, 18, -21, 7, -20, 26, -14, -3, -71, 1, 38, -26, -12, -4, 1),
    (11, 9, -3, -10, 22, -4, -11, 10, 32, -9, -2, -5, -1, 0, 21, 22, -24, 14, 1, 15, -27, 9, 12, -3, 16, 17, 10, 2, 6, -11, -14, -3, 12, -9, 13, 4, 3, -3, 5, 16, -19, 3, -9, 1, -22, 13, 1, -4, -11, 21, 2, -1, 11, -3, -4, 7, -9, -9, -1, 11, 12, 28, 0, 10, -10, -21, -4, 7, 0, 7, 13, -4, -9, -5, 5, 17, 7, 6, 28, 12, -8, -23, -2, 3, 15, -13, 19, 23, 12, -10, -6, -13, -4, -6, 17, -35, -13, 3, 3, 10, -3, 14, 1, 0, 1, -39, 2, 8, 19, 2, 4, 4, -13, -20, -40, 15, 20, 11, -4, -38, 14, 26, -12, 1, -16, 8, -8, 1, 18, -20, -6, 22, 14, 21, -7, -1, -20, -40, -42, 10, -4, -13, -1, -14, -40, -25, -7, 1, 7, 3, -16, -22, 2, 4, -21, 7, -10, -16, 6, 3, 5, 15, -31, -12, -7, 13, -15, 18, -41, -29, -10, -12, 12, -6, -1, -32, -10, -2, -12, 11, -4, -16, -11, 10, -13, 6, -53, -10, -8, 5, 1, 29, -24, -24, -10, -3, -13, -12, -17, -41, 11, -6, -20, 18, -13, -1, 6, 20, -14, -5, -55, -14, -12, -20, -24, 2, 0),
    (1, 28, -11, -5, -35, 5, 15, -21, -8, 17, 1, -1, 4, -29, -2, -13, -3, 7, 0, -22, 15, 0, -17, -19, 15, 27, 0, 23, -29, -11, -10, -20, -20, 7, -3, 4, 3, 4, -9, -16, 38, 23, 13, -12, -18, -2, 24, -25, 11, -5, 0, 24, -7, 10, 15, -2, -10, 7, -6, 10, 9, 23, -16, -2, 39, -5, 20, -24, -28, -5, -6, -11, -1, 12, 18, -5, -8, -23, -5, -18, 24, 2, -9, 13, -8, -6, 17, -3, -17, 16, -7, -15, 13, 10, -22, -21, -20, 24, -23, 5, -34, 0, 0, -6, -11, -16, -14, -23, 15, 12, 19, -2, 23, 5, 19, -20, 1, -4, -5, -31, -16, 27, -7, -19, -27, -11, 6, -20, 5, -5, -30, 18, 3, 31, 1, -10, 39, -33, 7, -22, -15, -2, -19, 5, -13, 15, -11, 15, 18, -2, 3, -16, 0, -14, 11, 17, 4, 18, -6, -4, -13, 26, 20, 11, -11, 17, -6, -13, -11, 14, -1, 3, -11, -5, 21, -17, 19, 5, -18, 2, -1, 4, 5, 4, -6, -10, 19, -18, -3, -5, -24, -2, -10, -7, -12, -9, -49, 5, 1, 4, 10, 14, -37, 7, -2, -4, 15, 6, 18, -19, 13, -16, -3, -11, 10, -6, 8),
    (-1, -20, 1, -21, -12, 16, -10, 7, -9, 0, 26, 14, 3, -14, -17, 21, 1, -3, 2, -18, 0, -4, -10, -1, -6, -40, 1, -2, -8, 28, 6, 16, -4, 2, 19, 1, -10, -19, -5, 35, 0, -26, 8, 2, 31, -6, 16, -8, -9, -18, -8, -9, 1, 20, 19, 23, -18, 1, 0, -1, 6, -25, -29, 22, 10, -28, 6, 12, 16, 16, 6, -3, 35, -6, -16, -17, -1, -15, -29, 1, 13, 17, -15, -8, -7, 36, -13, -24, -22, -11, 6, -18, -9, -17, -13, -7, 13, -38, -30, 3, -9, -19, -12, 34, 0, 21, 12, -13, -13, 17, -13, 0, -14, 1, -5, -9, 1, 9, 9, -2, 1, -22, -45, 13, -10, 6, 7, 30, -4, 9, 19, -12, -13, -7, -46, 6, -36, 7, 8, -7, -4, -12, 6, 15, 20, -12, -4, -26, -5, -14, -15, -2, 6, -7, -2, 5, 8, 14, 0, -2, -17, -52, 3, -6, 5, -8, -18, 14, -9, -22, -19, -6, -6, -9, -22, 8, -19, 14, -18, -6, 8, 29, -28, -7, -31, -17, 9, 9, -4, 10, -9, -5, -10, -16, -45, 11, -3, 9, 6, -7, -40, 1, 5, -16, 17, 13, -10, 7, -29, -21, 15, 0, 8, -23, -4, 14, -4),
    (-12, -4, 8, 6, 2, 0, -6, 29, -33, -5, 14, 14, -39, 1, -11, -1, 23, 12, -22, -9, -11, 12, 1, 14, 8, -5, -8, 2, 14, 6, -15, 12, -10, 24, 3, -6, -31, -20, -21, 4, 3, 2, -17, -7, -21, -3, 25, -3, 5, -18, -2, 3, -13, -6, -25, 21, -6, 9, 5, 14, -22, -12, 5, 9, -18, 12, -24, -3, 5, -7, 8, -10, 7, 4, 21, 10, -6, 2, 9, 7, -8, -5, 12, 5, -13, 2, -18, 6, 24, 8, 13, 4, 1, -4, -8, 3, -12, 9, 17, -2, 1, 23, -15, 9, -8, 15, 10, -4, -16, -27, -19, 15, 25, 8, 2, -6, 27, -4, 3, -7, -19, -13, 11, -2, -10, 13, 2, 14, -4, -6, 10, 7, 2, -24, -3, 5, 2, 13, 13, -17, -9, -2, 3, -4, 4, 6, 5, -4, 14, -7, -7, -2, -16, 9, 6, 2, 6, 1, -24, 2, 29, 14, 9, 18, -22, 10, 8, 15, -4, 23, -3, -18, 7, 13, -9, 8, -14, 0, -12, 5, -7, -14, -19, 18, 31, 6, 24, -13, 31, -27, 22, 0, -15, -2, 12, -9, 8, 11, 1, -2, 9, -1, 17, -1, -4, 6, 19, 7, 7, 0, 25, 16, 7, -2, 11, -10, -5),
    (-39, 0, -13, -50, -20, -15, 10, -30, 0, -3, -18, -39, 19, -32, -3, -12, -2, -4, -7, -14, 9, 2, -20, -2, -15, -28, -14, -16, 9, 10, 13, -23, -12, 24, 12, -25, 17, 0, 0, 1, 1, -22, -3, 8, 4, 3, 10, -26, -9, -1, -17, 17, 2, 7, 12, 3, -8, 7, 0, -5, 27, -5, -1, 12, -1, -36, 5, 23, -7, 15, 23, -5, -10, -3, -6, -46, -23, -10, -7, -24, 6, -5, 20, -22, 2, -8, -14, -3, -19, -6, 13, 7, 7, 2, -2, -24, 0, -10, -20, -15, 5, 7, 26, -26, -11, 39, 1, -41, 29, 10, 4, -25, 5, -11, 18, -8, 4, 9, 19, 10, -5, 0, -13, 15, 13, 3, 14, -2, -4, -8, 2, -2, 37, 28, 10, -19, 0, -14, 22, -7, -5, 7, -8, 20, 7, 0, 1, -18, -20, 17, -11, -27, 4, 31, -3, -25, -8, -4, 9, 7, -16, -22, 16, -30, -4, 13, 11, 6, 11, 7, -10, 24, 5, -4, 17, -13, -18, 19, 1, -13, 20, 16, 6, -26, -8, -18, 41, 13, -1, 9, -3, 12, 18, 4, -5, 12, -6, -16, -1, 4, 4, -14, 5, 7, 17, 33, 13, -9, -6, 8, 11, -8, -12, -5, -14, 4, -1),
    (-68, 28, 0, -48, -12, -21, -14, -38, 19, -32, -3, -5, -1, -67, 10, -10, -26, 11, -1, 7, 18, -24, -8, -10, -31, 40, -8, -37, -14, -1, -11, -27, -6, -27, -11, -15, -9, -59, -10, -24, -1, 14, 10, 6, 14, -1, -12, -9, -30, 24, -18, -34, -5, -23, -10, -37, -11, -5, -5, -21, 5, -20, 1, -2, -1, 22, 5, 9, 2, -5, -20, 17, -29, 13, -14, -10, -17, -9, 13, 4, 4, -9, 11, 7, -6, -6, 5, -5, -29, 21, -11, 10, -26, 2, -7, 6, -45, 48, -14, -36, 15, 2, -2, -5, 6, 15, 16, 2, 12, -2, -18, -16, -18, 32, 3, 9, -2, -13, -14, 14, -23, 44, -7, 1, 21, -13, -14, -14, -4, 4, -2, -24, 20, -5, -22, 17, -15, 24, 12, 5, 6, -1, 9, 8, -14, 7, 17, 17, 2, -12, 12, 22, 4, 9, 10, 18, -3, -13, 0, 22, 2, 34, -3, 11, -14, 17, 8, -2, -42, 34, 15, -12, 9, 6, -11, 23, 9, 0, 7, 2, 17, -9, -2, 12, 8, 43, -2, -14, 21, 9, 16, 2, -13, 28, 2, -9, 7, -9, 12, -14, 4, -12, 6, -13, 27, -2, 5, 18, -16, 18, -5, -4, 30, 21, 2, -3, 0),
    (15, 14, 3, 31, 21, 5, -4, 13, 11, -23, -2, -2, 12, -20, 1, 18, -3, -1, -16, 13, 10, 3, 8, -21, -3, 11, 10, 10, 17, 7, 5, -2, 4, -22, 4, 21, 6, -18, 13, 8, 16, 7, -16, 6, 23, 2, 12, -30, -1, 28, -4, -1, -19, -8, 2, -15, -15, 2, 1, 15, 4, -3, 1, 6, 11, 6, 9, -16, 24, 0, -14, -18, 0, 2, 24, 8, 14, -7, 17, 1, 7, 1, -10, 12, 24, -32, 31, 25, -7, 14, -12, 0, 18, 18, 2, -7, -13, 29, 13, -12, 6, 4, 17, -25, 20, -22, 1, 16, 21, -23, 24, 20, 14, 4, -38, -19, 46, -12, -16, 9, -4, 46, -4, -4, -2, -9, 16, -33, 22, -42, 0, -9, 7, 10, 14, -6, 2, -2, -32, -6, 22, -21, -15, -5, -23, 7, 5, -4, -6, 3, 24, 0, 0, 24, -22, 6, 22, -26, 13, 11, -1, 14, -1, -23, 0, -13, -10, 25, -28, 5, 22, -17, -27, -6, 6, -2, -11, 0, -26, 2, 28, -18, 10, 15, -7, 37, -38, -9, 13, -13, -1, 17, 3, 4, 12, -11, -2, -33, -15, -4, -16, -3, -3, 5, -4, 7, -8, 2, -9, 31, -53, 12, 9, -34, -12, 18, 6),
    (-38, 17, 15, -51, -18, -25, -5, -25, 5, 14, -26, -31, 30, -29, -17, 7, -3, -3, 0, -30, 12, -21, 6, -16, -15, 15, 0, -18, 11, 11, 17, -4, 13, -36, -20, -4, 38, -16, -15, -19, -14, -1, -7, -20, -11, -21, -18, -9, -12, 7, -1, 7, 14, 7, 3, -15, 20, -31, -21, -2, 7, -19, -8, -1, -5, -20, -3, -15, -12, -16, -15, -20, -30, -10, 18, 9, -4, 22, 19, -2, 25, 2, -29, -4, 9, -17, 14, -25, -17, 1, -16, -6, 20, -7, -23, -47, -10, -3, 25, 12, 3, 7, 29, 6, 40, -17, -17, 25, -6, -11, 30, -21, -13, 6, -14, -4, -5, 9, 7, -18, 4, 4, 26, 15, 0, 5, 3, 7, 31, -24, -17, 30, -10, 14, 35, -7, 8, 13, -12, 2, 9, 9, -25, -9, 25, 0, 5, 8, 2, 9, -4, 6, 10, -9, -14, 7, -10, -16, 18, 5, 7, -10, -3, 2, -8, -5, 0, -19, 29, 3, 9, 16, 19, -6, -15, 17, -2, -14, 11, 13, 4, 17, 27, -8, 1, 16, -9, 19, -8, 8, -13, 4, 8, 8, 4, 10, 8, 14, -17, 33, 2, -8, 4, 9, 9, 9, 20, 14, 12, 16, -8, 14, -14, 3, 14, -15, 5),
    (-20, -3, -5, -4, 12, 8, -1, 1, 16, 7, 18, 0, 9, -2, 11, 14, -18, 7, -4, 19, 2, -2, 10, 19, -38, -18, -25, -6, 6, -9, -27, -27, 8, -5, 21, -36, 9, 1, -8, -30, -21, 8, -15, 9, 9, 3, -1, 27, -30, 6, -30, 2, -9, 0, -21, -19, -18, -14, 9, -36, 3, -13, -18, -12, 1, -10, 0, -28, 25, -26, -8, 19, -23, 8, 20, -9, 4, 1, -9, 12, 10, 17, 12, -10, 3, 19, 21, -7, 5, 18, -1, -15, 31, 3, -5, 34, -34, 22, -12, -16, 21, -14, -16, -6, 8, 2, 17, -41, 31, -3, -13, -8, -1, -1, -14, -6, 31, 16, 5, 26, -18, -6, -22, 14, -9, -17, -18, -19, -16, -13, 6, -10, -7, 6, -39, -23, -3, 3, -18, -9, 5, -11, -8, 5, -5, 22, 0, 2, -6, -6, 2, 8, 7, 18, 18, -3, -13, -1, -2, -13, 9, 9, 15, 0, 11, 15, -3, 31, -23, 19, -19, -14, 2, -23, 5, 5, 10, 14, 7, -24, 39, -8, 0, 7, -2, 12, 12, -6, 29, 16, -5, 30, -8, -23, -22, 17, -16, -14, -13, -10, -6, -21, -24, 0, -2, 2, -6, -17, -7, 26, -51, -18, -1, -3, 6, -1, 0),
    (-25, 11, -16, -4, -5, -3, -43, -19, 25, 26, -21, -53, -44, -23, 18, -10, -16, -31, -10, -23, -25, -9, -21, -6, -2, -9, -11, 5, 10, -6, -13, -10, 1, -1, -19, -37, -43, -12, 14, -9, 3, 1, 3, -13, -42, -28, -12, -5, 2, 25, 3, -3, 8, -32, -20, -39, -2, 8, -15, -49, -25, -4, -17, -35, -26, 1, -4, -6, -55, -19, -1, 4, 35, -2, 11, 22, -6, 2, -27, 25, -6, -7, 17, -30, -31, -18, 10, 8, -14, -14, -8, -2, 0, -1, 14, -25, 43, 14, -14, 27, -6, 7, -26, 24, -26, 26, 5, -8, -45, -23, -13, -1, 14, -9, 12, 13, -12, -18, -7, -38, 34, 0, 1, 23, 2, -30, -32, 7, -21, 21, -11, -4, -43, -5, -27, 11, 8, -4, 16, 16, -17, 6, -11, -40, 24, -7, 11, 23, 6, -4, 16, 18, 14, 8, 6, -16, -12, -9, 1, 26, -5, 9, 7, 7, -31, 2, 12, -14, 27, 19, 13, 28, 2, 13, 21, -3, -4, 6, -17, 1, -4, -28, -3, 49, -2, 10, 8, 15, -17, 13, 4, -9, 8, 6, -4, 15, -2, 8, 5, -5, -10, 12, 11, -3, -2, -7, 3, 13, -5, -7, 15, -10, -22, 14, 6, -1, -1),
    (12, -15, 6, -6, -5, -26, -13, 1, 3, -20, 14, -8, -3, 25, -16, -14, -10, -14, 4, -9, 33, 5, 1, 3, 5, 12, 17, 6, -8, -26, -14, -14, 10, -4, -5, 37, -3, -13, 7, -31, -5, -2, -7, -16, -6, 9, -2, 0, -1, 20, 31, 3, 20, -7, -1, -19, 11, -40, -28, 21, 11, 15, 22, -12, 11, -4, -3, -9, 0, 4, 3, -16, -23, -1, -16, 0, -15, -10, -17, 14, 14, 9, 6, -9, -9, 16, -3, 7, -16, 4, -14, -18, -9, -7, -19, 0, -9, -10, 16, -9, -15, 7, -6, 1, 27, -6, -26, 14, 8, -13, 16, -6, -1, -2, 7, -19, -2, 1, -12, 10, -25, 1, 23, 3, -15, -4, 14, 12, 24, -47, -23, 30, 14, -8, 42, 1, 6, 8, 12, 10, -2, -10, -6, -1, -7, -20, -1, -16, 3, -3, -13, -13, 3, 15, -14, 9, -5, -6, 2, 0, -9, -18, 5, -31, 16, 8, 6, -21, -20, -16, 8, 12, 8, 5, 19, 5, 23, -2, -11, 15, 8, 18, 4, -11, 9, 8, 16, -22, 0, -13, -5, -10, -22, -13, 26, 12, 22, 20, 21, 4, 20, 0, -7, 13, 6, -9, 37, -1, 2, 8, 3, 5, -6, 2, -11, 25, 0),
    (-8, -20, 7, 8, -12, 30, -10, 20, 12, -17, 18, 19, -6, -4, 25, 1, -8, -7, -21, 13, 19, 9, -2, 0, -17, -21, 1, -4, 8, 22, -13, -3, 14, -23, 21, 0, -1, -18, -8, 13, -7, -2, -4, 7, 17, 10, 22, 13, 3, -13, -37, 7, 0, -12, -15, -21, -19, -11, -1, -6, 8, -9, -33, 13, -14, -13, 15, 7, 39, 3, 25, -5, -2, -14, 13, -19, -5, -1, 4, 6, 17, 1, 7, 31, 7, -1, 13, -1, 1, -33, -7, 14, 7, 7, 0, -6, -39, -24, 11, -37, 15, 7, -20, 0, 38, -8, 17, 13, 4, 0, 14, -14, 3, -9, -7, -5, 28, -6, 6, 35, -12, -41, -19, -3, 4, 12, -18, -18, 7, 7, 15, -24, 0, -7, -21, 10, -1, -33, -8, 17, 52, -1, 23, 14, 0, -14, 17, -11, -23, -5, 5, -4, 4, 3, 15, 21, -9, 1, 9, -6, -1, -20, -15, 4, 6, 1, -1, -36, -23, -19, -4, -20, 2, -2, -4, 8, -2, 2, 17, 8, -1, 14, 16, -9, 9, -24, -20, -11, 23, 10, -10, 15, -17, -30, -15, 3, -3, 15, -17, 11, 0, 7, 21, -19, -9, -9, -10, 15, -12, -11, -9, 16, -2, 0, 23, 5, -6),
    (-8, -9, -22, 0, -4, -16, -13, -9, -26, -10, 8, -30, -1, 13, -17, -16, 19, -17, 11, 18, -20, 13, 1, -2, 16, -23, -23, 17, 4, -14, -18, -8, -20, 4, 22, 1, -15, 1, -34, 8, 23, -36, 14, 4, -17, 0, 14, -12, 16, -9, -4, 5, -6, 5, 4, 1, -7, -4, 10, 20, -17, -18, 5, 5, 19, -21, -33, -7, 9, -8, -7, -15, -5, -13, -31, 6, 20, 10, 1, -4, -35, -21, 1, -33, -6, -15, -38, 1, -6, -32, 4, 20, 20, 17, 24, -11, 5, -20, -28, 9, 8, 6, -8, -5, -8, -13, 14, -5, 4, -27, -32, 42, 29, -42, 8, -3, 23, 21, 29, -34, 3, -14, -5, 8, 9, -9, -3, -24, -4, -11, -2, 18, 3, -4, 12, 12, 22, -30, -15, -5, 23, 9, 6, -28, -16, -9, 0, 5, -9, 7, 4, -12, -30, -10, 4, -14, 4, 1, -16, -14, -14, -12, 10, -7, 15, 10, 13, 14, -27, 16, -4, 1, 12, 32, 16, -23, -7, -24, 13, -2, 36, -16, -2, 9, 5, -4, 6, -10, 31, -5, -5, -18, -18, -26, 9, -8, -3, -7, 1, -20, 16, -17, -24, -2, 8, 18, 15, -1, -5, -11, -44, 8, 3, -19, -21, -25, 0),
    (-25, 28, 38, -36, -10, -13, -20, -23, 13, 19, -15, -21, -5, -8, 8, -31, -7, 8, 0, -14, -30, 0, -13, 20, -13, 27, 1, -2, -1, -19, -8, -13, -4, 16, 4, -28, -14, 22, 5, -41, -17, 2, 15, 3, -47, -3, 1, 40, -9, 11, -5, 0, -8, -11, -6, -7, 7, 16, 0, -17, -9, 8, 4, -31, -19, -5, 11, 5, -36, 19, 7, 7, -15, 30, -1, -25, -14, 0, -26, -9, 0, 29, -11, -31, 17, 10, -2, -25, -20, 6, 22, -7, -33, -15, 9, 2, 6, 27, -9, 25, 6, -3, -19, 6, -4, 28, 21, -31, -13, -7, 7, -15, -27, 26, 21, -4, -53, -16, -2, -2, 7, 14, 1, 15, 5, -3, -28, 28, -11, 6, -4, -26, -12, -8, -4, -4, -13, 6, 11, -1, -29, 17, 25, -5, 25, 16, -11, 2, 4, -3, -20, 16, -17, 12, 11, -12, -4, -1, -7, -5, -25, 6, 20, 2, -10, -11, 15, 5, 23, 18, -10, 21, 13, -3, -30, 22, -24, 22, -9, -16, -2, -18, -4, 2, -27, 13, 22, 17, -22, 9, 25, 1, 4, -5, 1, 14, 19, 1, -4, 24, -15, 4, 18, -6, 8, -13, -5, 18, 1, 0, 18, -2, 4, -7, 7, -2, 4),
    (30, 8, -7, -7, -16, -26, -8, -21, 7, 17, -22, -7, -10, 51, 1, -16, -23, -15, -11, -5, 9, 1, -2, -41, 29, -30, -5, 8, 16, -13, 9, -19, -15, 15, -6, -13, -19, 30, -8, -13, 42, -23, 3, -9, -27, -3, 1, -33, 23, -5, 23, 9, -12, -17, 20, -14, -15, 16, 1, 8, -17, -7, -10, 3, 30, -2, 24, -1, -30, 8, -1, -3, -3, -19, -19, -11, -6, 2, 0, 11, -18, 15, 19, -50, 7, 14, -6, -4, -10, -7, 3, -2, -30, 18, 3, -11, -7, -47, -21, 1, -13, -7, 14, -10, 6, 10, 1, -23, 4, -11, -17, 8, 29, -7, 0, 25, -30, 6, 22, -15, -10, 8, -9, -20, -10, 10, 13, 1, -7, 16, 17, 1, 0, 1, 17, 15, 25, -13, -2, -4, -18, 13, 8, 0, -19, 7, -8, 9, 9, -3, -3, 6, -22, 3, 17, -3, -6, -18, -15, -25, 13, -5, 6, 8, -9, 16, 9, -2, -5, 8, -20, 7, 4, -5, 15, 3, -24, -19, 9, 4, -6, 7, -7, 7, 13, -29, 6, 3, -16, 10, 5, -13, 13, 8, 14, -4, -2, 1, 11, -9, 3, -19, 19, -2, -9, 7, -1, 0, -5, -25, -3, -9, -2, -1, 5, 4, -4),
    (-14, 7, 16, 1, 12, 19, 27, 3, -20, -13, -13, 16, 14, -3, 13, 11, 0, -23, -17, 7, 16, 16, 22, -13, -5, 27, -4, 13, -8, 6, 23, 4, -8, -46, -11, 6, 26, 16, 16, 11, -12, -17, -34, -2, 11, 9, 6, -25, 32, 27, -3, -2, -25, 2, 1, -4, 4, -45, -10, 5, 5, 12, 0, -5, -6, -28, -39, -3, 12, -5, -9, -19, -59, -16, -8, 3, -9, -9, 2, -37, 0, 8, 6, -10, -7, -25, 2, 4, 6, 8, -30, -1, 27, 27, -10, 26, -50, 1, -9, 2, 13, -16, 22, -30, -11, -13, 6, 6, -2, -17, -12, 10, -16, 12, -49, -20, -5, -5, 10, 11, -24, -18, 21, 5, 2, -15, -3, -26, -31, -27, -9, 3, -27, -9, -29, -7, 12, 40, -40, -17, -17, -11, -21, -6, 11, 0, 21, -22, -15, -14, -7, -2, -11, 9, 4, 7, -35, 25, -2, -24, -7, 7, -4, -3, -3, 26, -11, 8, 9, -2, -15, -43, -7, 9, -13, -3, -17, 12, 1, -6, -31, 32, -3, -27, 3, 3, -5, 2, -2, 10, -2, 19, -17, -8, 7, -5, -8, -20, -19, 8, -15, 2, 21, -46, -7, 3, -38, 4, 18, 5, -12, 13, 0, 22, -4, 0, 0),
    (-6, -12, 0, 1, -5, 15, 7, -15, 7, 5, 11, -12, 14, -7, 13, -3, 6, 9, 4, 1, 13, -6, 16, 27, -29, -7, -17, -8, 21, -1, 23, -18, -22, 36, -1, -20, 26, 15, -3, -4, 5, 16, 12, -9, 0, -17, -8, 22, -6, 5, 19, 5, -10, 3, 4, -4, -25, 3, -14, 16, 5, -2, 1, 11, -3, 22, -17, -2, 14, -5, -20, -6, 26, 2, 16, 18, 7, -7, -3, -4, 10, -23, -20, 23, -3, 25, 24, -19, 0, 10, 8, -12, -34, -4, 17, -13, 12, 14, 16, -23, -6, -13, -10, 17, -3, 20, 18, -6, 15, 40, -17, -22, -14, 17, 15, 6, -29, -24, -20, 29, -26, -13, -7, -12, 24, 8, -27, -9, 4, -3, 13, -3, 5, 21, -13, -17, -8, 32, 5, -17, 9, -9, 12, 16, 10, -11, 19, 20, -6, -5, 5, 3, 3, -11, -4, 17, -24, 5, 13, -7, -10, -7, -19, 3, -37, 0, 5, -29, 36, -24, 13, -23, -9, -19, -17, 27, -13, -18, 13, 31, -29, 23, -28, 1, -14, -18, -8, -5, -39, -25, -18, -6, 19, 8, 3, 5, -20, -14, -41, 1, -35, 8, -11, -4, -28, 16, -28, 4, -17, -2, -48, 7, 3, 2, 6, 5, -8),
    (27, 5, 11, -15, -11, -9, -19, -1, 14, 32, -11, 6, -5, 26, -6, -22, -4, -1, 15, -12, 6, -3, -18, -1, 25, 2, -21, 7, 0, -12, -25, 23, 13, 17, -21, 5, -6, 7, 4, -7, -5, 17, 8, -15, 6, -7, -11, 6, 14, -3, -34, 6, 12, -7, -21, 26, 15, 4, 1, 18, -2, 5, 5, 2, -13, 16, 18, 7, -16, -24, 5, 2, 28, 21, -35, -4, 15, 0, -27, 21, -18, 30, -4, 0, 3, 32, -31, 15, -14, -4, 32, 16, -2, -24, -3, -2, 27, 43, -17, 6, 9, -5, -24, 12, -21, 28, 3, 22, 6, 28, -14, -4, -5, 19, 37, -6, -14, -7, -14, 5, 12, 30, -25, 7, 9, -22, -21, 4, 0, 9, -12, 32, -8, 23, 8, 0, -20, 29, 15, -24, 2, 6, 4, -6, 19, 5, -37, 7, 8, -14, -15, -3, -12, 13, 1, 0, -19, -1, -18, -6, 5, -3, 14, 23, 13, 24, 26, -3, 22, 46, -28, 17, 6, -8, -24, -15, -22, 17, 15, 1, -20, 0, -19, 6, -21, -3, 31, 12, -2, -19, 17, -2, -6, 23, -25, 17, 0, -6, -20, -3, -18, -1, 10, 12, 9, 18, -7, 11, 0, 19, 2, 6, 3, -2, -4, -13, -16),
    (7, 1, 20, 1, -13, -2, 7, -6, 5, 7, -17, 5, -5, 37, 15, -16, 12, -17, -11, 8, 11, 6, 2, -35, 23, 6, 3, 12, -4, 3, -13, -1, 12, 14, 11, 4, -4, 39, 25, -25, -8, -4, -1, 18, -11, -24, 11, -26, 6, 25, -3, 12, 9, 5, 14, 22, 5, -2, 8, 7, -3, -5, 9, -25, 5, -27, -13, -8, -9, -17, 17, -16, 41, 14, -2, 12, -18, -11, -16, 1, -9, 8, -13, 9, -19, 41, 16, -39, -4, -10, 10, -6, -16, -13, 22, -63, 35, 18, -11, 5, -5, 12, -18, 21, -11, 21, 2, -1, -34, 34, 13, -37, -18, -2, 5, 18, -43, -15, -15, -18, 25, 12, -5, 26, 0, -7, -23, 25, -23, -7, 16, 0, -26, -9, -24, -20, 10, 0, -61, -1, -25, -9, -13, -6, 15, 36, 14, 3, -5, -14, -11, 20, -23, -6, -4, 10, -26, 26, -15, 0, -26, -60, 12, 16, -22, 18, 4, -25, 18, 23, -29, 3, 1, 12, -16, 17, -7, 6, 26, -3, 11, 18, -22, 3, 1, -36, 19, -12, -18, -12, 12, -11, 6, 10, -37, -1, 8, -7, 9, -4, -18, 23, -16, -11, -16, 10, -21, -4, -6, -26, -53, -6, -8, -5, -27, 10, 0),
    (-10, 3, 7, -2, -3, -4, 2, -9, -4, -12, -16, -7, 10, -29, -2, -12, -7, -7, -21, 1, -25, 18, 13, -13, -9, 6, -15, -17, 8, 0, 26, -18, 2, -31, 6, -9, 23, -24, 3, -28, -35, -20, 0, -3, 1, -4, 2, 2, -1, -10, -13, 10, 24, 33, 26, -25, -1, -29, -24, -17, 18, -15, 14, 4, -3, -11, 3, 1, -9, 0, -2, 3, -6, -1, 7, -3, 6, 38, 5, -7, -5, -7, -21, -13, 17, -27, -1, -14, -5, -5, -7, -8, -2, 15, -11, -19, -2, 1, 4, 6, 6, 23, 11, -10, -1, -32, -5, -1, 6, 1, 7, -41, -38, -4, -8, 15, -9, 2, 0, 14, 4, -12, -10, 15, 9, 33, 28, -10, -3, -26, 3, -10, -9, 0, 26, -16, -22, -26, 1, -13, -24, -5, 26, 5, 18, 22, -5, 6, 12, 8, 13, -9, -24, -17, -14, 3, -6, 17, -11, -9, -20, -6, 3, 18, -8, 15, -4, 29, 4, 11, 2, 10, 11, 4, 2, 6, 0, -18, -8, -4, -3, 0, 4, -10, -27, -7, 2, 8, -19, 18, 6, 8, -2, -14, 0, 3, 1, 29, 16, -4, -10, 11, -11, -12, 6, -11, 13, 1, -9, -2, 14, 2, -15, 6, 23, 21, -1),
    (10, 0, 20, 16, 0, -13, 9, 18, 5, -1, -2, 10, -6, 9, 6, -4, -8, -19, 18, 21, -35, 22, 9, 7, 3, -10, 5, 12, 7, 10, 0, 2, 2, -16, -12, 21, 14, -6, 11, 10, 18, -5, -11, 18, 13, 10, 2, 10, -7, 19, -9, -2, -12, -19, -10, 7, 4, 8, 13, 9, 1, 6, 8, -14, -5, 49, -5, 1, 16, -22, -16, -2, 1, 4, 9, 20, -5, 8, 12, -1, 2, -15, 3, 18, 7, -4, 2, -14, 1, 14, 16, 6, -17, 4, 23, 29, -11, 9, -6, 9, 12, -3, 29, -17, 23, -21, -37, 10, -1, -13, 37, 0, 3, 1, -14, -14, -4, -3, 5, 7, 2, 41, 1, -18, -15, -28, -6, -11, 1, 14, -7, 2, -12, 14, -3, 2, -6, 38, -20, -26, 9, -13, -19, -2, -10, 0, 0, 11, 20, -3, 14, 4, 3, -9, -10, 13, -5, -28, 4, -1, 16, 8, 4, -3, 12, 16, 25, 26, -3, 6, 10, 8, -2, 3, 8, -15, 6, -27, -11, 9, -30, -20, 29, -23, 10, 6, -21, -20, 5, -1, -4, 11, 6, 30, 2, -20, -17, -23, 9, -14, -9, 9, -23, 2, 1, 12, -1, -2, -7, 24, -30, -9, 22, -22, -2, -4, 2),
    (-43, 38, 8, -25, 0, -7, -12, 5, 1, 4, 8, -10, -2, -33, 16, 10, -27, -7, -16, -21, 6, -16, -22, -25, -12, 36, -3, -10, 11, -15, -10, -4, 0, 10, -8, 16, -31, -30, 30, 15, 15, 36, -26, -19, 7, -3, -11, -2, -4, -2, 23, -5, 11, 11, -10, 2, 1, -2, -21, 6, -18, -8, -1, 6, -12, -11, -8, -11, 0, -2, -6, 7, -27, 36, 4, 10, 1, 6, 0, -13, 18, -4, -27, 18, 18, -12, -19, -16, -7, -7, 6, -6, 6, -24, 3, 0, 9, 6, -18, -10, -1, 13, 4, -13, -18, 13, -18, 15, -29, 21, 3, 1, -2, -18, 15, -8, 21, -15, -11, 5, 17, -53, 9, 1, -8, -4, -38, 5, -1, -25, 3, 8, -4, 0, -8, 6, -8, -37, 11, 13, -11, 6, -12, -14, -42, 4, -19, 3, 21, 13, 32, -8, 0, 13, -22, 15, 5, -9, 13, -13, -22, 32, -12, -8, 13, 6, -21, 8, -30, 7, 6, 3, 24, 21, 14, 3, -7, -31, -30, -20, 26, -19, -18, -6, -16, -7, 19, 4, -16, 4, -3, 9, -3, -9, 1, 24, 27, 14, -31, 4, -10, -17, 27, 1, 25, -20, -13, -20, -22, -46, 3, 7, -28, 10, -9, -17, 4),
    (11, -24, 12, -7, 8, 17, 15, 16, 14, 4, 8, 16, -22, -8, 16, 2, 17, -26, -23, 3, -5, -11, -6, 5, -14, -8, 0, -17, 11, -3, 18, -4, 8, 7, -1, -12, -10, -13, 5, 9, 11, -33, -31, 4, 22, 16, 22, -7, -7, 5, -24, -13, 6, -11, 5, -26, -6, 25, -6, -20, -9, 3, -21, 15, 13, -13, -18, -2, 30, -4, 4, 0, 3, -25, 5, -8, -25, -16, -4, 23, -3, 20, 21, 11, -15, -12, -1, -5, 30, -71, -6, 17, 8, 9, -14, -25, -23, -34, 6, -21, -2, 13, 5, 8, 19, 33, 9, -4, -32, -25, 20, 18, 33, -9, -15, 6, 39, -4, 7, -8, -33, -14, -11, -22, -7, 16, 8, -8, 12, 30, 17, -23, -36, -18, -6, 22, 19, -5, -1, 5, 46, 21, 14, 7, 3, -13, -11, 3, -8, -23, 3, 0, -5, 16, 13, 0, -2, 4, -21, -3, 8, -12, 28, -7, 5, -13, -6, -54, 17, -18, 9, 6, -20, 3, -15, 6, 8, 29, -6, -1, -33, -5, 8, -5, 22, -24, 20, 1, -16, 6, 5, -29, -3, 6, 23, -1, 1, -11, -2, -3, 0, 21, 10, -13, -5, -1, 9, -5, 12, -28, 22, -8, 1, 8, 3, -4, -3),
    (25, 14, 3, -5, -9, -7, 0, -18, -16, 7, 17, -4, 27, 15, -6, -20, -1, -27, 12, -26, -30, -10, -5, -18, -1, 35, -15, -2, -1, -11, 14, -23, -34, -10, 25, -16, 34, 20, -18, -6, 7, -30, 31, 17, -19, 17, 10, -22, -3, 27, -26, 2, 17, -7, -9, -22, -11, -13, -5, -6, 25, 19, -6, -10, 10, -15, 28, -14, 11, 13, -8, -22, -8, 35, 0, -21, -29, 5, 31, -36, -9, -10, 17, 19, 29, 2, -2, -9, 19, 11, -4, -9, 16, -10, 9, -8, -22, 40, -16, -28, 8, 14, 27, -38, -17, -22, 19, 6, 31, 31, -12, -21, 8, -22, 17, 4, 28, -8, 23, 6, -6, -1, 7, -13, 15, -16, 3, -24, -9, -2, -5, 0, 17, 30, -3, -14, 1, -24, 4, -4, 21, 3, 18, -3, -2, 16, -4, -19, -21, -4, 29, -10, -20, -14, 2, 15, -10, 8, 8, -3, -2, -24, -11, -3, 3, 6, -14, -30, 4, -2, 1, -15, -16, 15, 12, -28, -29, 6, -14, -3, -4, 28, -11, -27, -3, -37, -14, -1, 6, 13, 6, 14, 11, -28, 15, -5, -14, -13, -4, 4, -12, 7, -20, 4, -2, 8, 3, -8, -9, -27, 1, 6, -23, 1, 10, 11, -3),
    (-3, 27, 12, 11, 5, -13, 14, 2, -20, 21, 13, 1, -9, 21, -31, 13, 37, -18, 1, 3, -7, 5, 4, 12, 3, 26, 9, -14, -12, -17, -1, -15, -20, 7, 18, 21, 8, 40, -29, -2, 12, -3, 23, 2, 1, 13, 2, 8, -8, 9, 5, -15, -4, -5, -9, -6, -20, 11, 1, 28, 21, 37, -18, 9, 8, -14, 18, -15, 25, -2, 5, 20, 1, 16, 9, 3, -5, 16, 9, -9, 10, -21, 3, 19, 7, 9, 0, -5, 22, 11, 1, 12, 4, -5, 21, -22, 0, 28, 31, -12, -16, -5, 9, -33, -6, -9, 15, 22, -2, 4, -9, 10, 7, 22, 2, 20, 9, -10, -1, -10, 4, 11, 17, -6, -19, 1, 3, -7, -6, -20, 18, 27, 10, 19, -3, -17, 10, 11, 3, 11, 17, 0, 12, 7, -20, -20, 19, 7, 6, -1, 26, -6, 4, 7, -28, 4, -4, -15, 6, -15, 22, 10, -18, 8, -26, 8, -1, -9, -7, -9, 7, -28, -12, 15, 10, -24, 20, -31, 7, 25, 5, 1, 7, -25, -5, 0, -22, 14, -12, -16, -14, 13, -1, -19, 21, -3, -7, -1, 21, -2, 25, -24, 10, 10, 1, -12, 12, -3, -4, -9, -22, 17, -3, 9, 4, -11, -5),
    (-2, 32, -19, -14, 4, 12, 9, -28, -6, -3, -8, -39, 26, 17, -5, 14, 12, 5, 2, -17, 45, -19, -8, -24, 32, 29, -27, -10, -18, -8, 10, -14, -8, 2, -17, -57, 2, 33, -4, -1, 9, -4, -9, -2, 44, -16, 13, -27, 29, 7, -7, 3, -14, -8, 19, -1, -6, -11, -1, -28, -14, 7, -12, 0, 22, -13, -12, 7, 6, 9, 15, -36, 26, 2, -14, 0, -4, 1, 5, -7, -42, -13, 13, -47, -2, 20, -18, -10, -6, -28, 5, 11, 11, -11, 22, 4, 31, -4, -54, 6, -7, -6, 16, -20, -33, -3, 18, -36, -14, 26, -29, -1, 15, -21, 26, 4, -11, 13, -3, 1, 21, 5, -24, 13, 4, 9, 24, -8, -15, -5, -9, -8, -1, -1, -11, 6, 9, -4, 19, -1, -12, 16, 6, -9, -3, 9, -10, -3, 4, 3, 11, -9, -7, 0, 6, -22, 0, -2, -23, 9, -1, 3, 1, 9, 9, 1, -1, 19, 7, 4, -20, -2, 13, -12, -7, -16, -20, 4, -1, -20, 11, -11, -31, 3, 8, 5, 16, 12, 12, 14, 16, 12, -11, 4, -20, -1, 4, 14, 21, -12, -7, 14, 21, -9, 7, -11, -13, -3, 4, -1, 26, -9, 7, 7, 18, 20, -2),
    (-12, 24, 17, -7, -15, -1, -11, -13, -2, 14, -6, 18, -1, -22, 3, -12, -6, 10, 6, -27, 13, -18, -16, -15, 1, 27, 31, 1, -11, -6, -12, -6, 13, -14, -16, 37, 12, -2, 22, -14, 18, 18, 2, 8, 7, -14, 5, -20, 1, 15, 18, -14, -7, 15, 7, 11, 6, -12, 10, 19, 5, 5, 16, -4, 13, 12, -3, 15, -6, -10, -13, -8, -15, 16, 25, -23, 9, -13, 10, 10, 19, 19, -12, 19, 13, -20, -2, -7, -13, 3, 7, -6, -9, -19, -26, 0, -21, 38, 29, -15, -13, 11, 15, -11, 33, -13, 1, 61, 4, 0, 40, -35, 5, 26, 18, -13, -22, -8, -5, 5, -1, 29, 26, -17, 6, 4, 2, -14, 6, -12, -16, 27, 4, 0, 20, -27, -7, -3, 19, 7, -22, 11, 7, 3, -7, 24, -7, -11, -8, -5, -11, 3, 11, 3, -13, 9, 27, -16, -9, -9, 1, 16, 29, -16, 5, 6, 14, 4, -25, 23, 20, -13, 9, 18, 3, -19, 6, -9, -5, 19, 9, 8, 27, -9, -13, 16, 17, 5, -11, -8, -20, 13, -7, 5, 4, -6, -10, -14, -2, -11, 0, -12, 9, 17, -3, 18, 1, -23, -12, -5, 16, 8, -6, 18, 10, 4, -3),
    (-43, 10, -36, -42, -21, 11, -8, -12, -15, -13, 10, -35, -1, 2, -20, -19, -21, 22, 1, -7, -2, 8, 6, -25, 0, -49, -27, 13, -9, -28, -34, -4, -34, -2, 7, -30, -16, 4, -26, -30, -10, -33, 4, 8, -52, 4, -2, 2, 16, -26, -6, 34, -17, -4, -6, 4, -15, 3, -2, -5, -24, -15, -10, -26, 15, -32, -11, 28, -25, 26, -4, -20, -24, -39, -41, -1, -2, -17, 17, 0, 29, 1, -18, -37, 12, 17, -2, 4, -23, 4, 7, -21, 4, -14, -9, -29, -3, -48, -34, 18, 17, 6, -1, 8, 2, -23, 16, -70, -5, 0, -27, 27, -18, 3, -3, -10, 6, -2, 18, -18, 0, -31, -12, 0, 14, -8, 15, -12, -20, -1, 9, -23, 5, -18, -24, 29, 19, -45, -2, 11, 2, -4, -2, -40, 6, -48, -3, 14, -8, 9, 17, 9, 7, -11, 12, -5, 8, -8, 20, 25, 0, -10, -22, -5, 36, 1, 2, 1, -17, -44, -4, 13, -5, -7, 19, -8, 10, -27, 11, -24, 20, -26, 1, 25, -13, 10, -3, 6, 34, 13, -9, 8, -27, -9, -10, -6, 25, 8, 0, -15, 5, -5, 19, -5, 30, -9, -9, 18, 7, 8, 2, -1, 30, 11, -4, -5, -1),
    (-10, 8, -13, 2, 0, -17, 13, -30, 25, -15, -17, -2, -5, -67, 27, 11, -8, 20, -8, 8, 26, -26, -11, -5, -2, -11, -19, 3, 4, 8, -18, -24, 19, -31, -8, 21, -5, -42, 25, 16, 5, 5, -12, 11, 32, -2, -1, -7, 10, 17, -12, 2, 10, -40, -1, -8, -10, 8, -26, -15, -23, 26, 13, 13, -19, 5, -20, -29, -9, -15, -28, -28, -5, -31, 6, 10, 19, 12, 16, -1, 22, -7, -6, -29, -17, -31, 36, 19, -19, -3, -23, 7, 6, 9, 15, 8, -30, -32, 6, -9, 14, 20, 7, -8, 29, -15, 4, 13, 22, -18, 18, 30, -1, 13, -31, -11, 29, 15, -9, 8, -23, 2, -8, -23, 17, 4, -7, -34, 8, -7, -9, -6, 19, 3, 28, 25, 3, 32, -23, -23, 3, -12, 10, 5, -17, -12, -5, -14, -5, 4, -7, 0, -16, 15, 13, -7, -15, -8, -9, -4, 9, 2, 3, -15, -6, 8, -10, 19, -12, -5, -1, -21, -18, 4, 6, -7, -10, 17, -7, 7, -11, -3, 12, 16, 5, 7, -20, 12, 11, -6, 15, 25, -21, 7, -2, -31, 11, -10, 9, -13, -10, -7, -13, 2, 18, -5, 18, 7, 1, 17, 0, -26, 55, 12, -5, 20, 5),
    (-23, -23, -2, -19, 11, -8, -8, -8, 12, -17, -7, -8, -12, -43, -4, -11, -16, -17, -4, 9, 8, 8, -9, -39, -14, 10, -2, -12, -9, 16, 24, -31, 17, -3, -15, 6, 20, -42, 15, 15, 21, -12, 7, -2, 12, 18, -9, -29, -9, 21, 8, -8, -7, 13, 4, -9, 6, -26, -3, 16, 30, -30, 7, 17, 2, 4, 20, 7, 8, 0, -9, -29, -20, 6, -26, -25, -2, 24, 18, -11, -6, -26, -22, -3, 15, -24, -9, -13, 0, -19, 9, -10, 23, 11, 19, -24, -30, 32, -1, -7, 3, 28, 29, -29, 21, -18, -18, -7, 36, -3, 26, 3, 17, -14, 5, 6, 7, -14, -9, 3, -25, 40, 0, -8, -5, 21, 2, -4, -14, 1, -15, 3, 21, 20, 16, -24, 6, -1, 4, -12, 12, -8, 16, -7, -11, -3, -18, 1, 17, 13, 30, -5, -3, -14, -6, 1, 14, -16, 5, -4, 13, -7, 1, 16, -2, 2, 9, 2, -22, 16, -6, 2, 15, 23, 15, -16, 3, -27, -4, 0, 17, 1, 27, -15, 3, -5, 10, -13, 3, -9, 17, 10, -17, 29, 3, -13, 6, 11, -6, 7, -21, 11, 5, -7, -2, 21, -29, -15, 7, -16, 8, 11, 15, -4, -13, 15, -2),
    (-10, -38, -3, -3, 17, 5, -1, 3, -4, 6, 29, -1, -21, -28, -11, 15, 6, 0, 4, 5, 20, 6, 5, 5, 0, -14, -9, 14, 17, 9, 5, -2, 12, 8, 10, -3, -6, -55, 11, 26, -2, -10, 4, 19, 20, 20, 10, 7, -10, 13, 7, 13, 20, 21, 0, -5, 11, -2, 18, 0, 10, -14, 17, 18, 0, -20, 5, 7, 23, 22, -11, 3, -14, -41, 6, -5, -3, 6, -28, 7, -13, 29, 11, -4, 13, -8, -14, 9, -16, 2, 1, -6, 20, -9, -26, -24, -24, -37, 0, -14, -2, 22, 2, -2, 13, 4, 22, -5, 10, -18, -34, 24, -21, 0, 2, 2, 43, 12, 8, 2, -11, -12, -3, -14, 13, 1, 6, -9, 6, 2, 2, 4, 8, -4, -20, 13, -2, -31, -11, -7, 29, 6, -6, 6, -1, -1, 14, 1, -18, -9, -22, 15, 24, 25, -6, 1, 13, 33, 16, -37, -13, -17, 5, -37, 7, -28, -3, 10, 11, -23, -4, -16, -14, -8, -14, -4, 5, 6, -22, -1, 16, 24, -12, -6, -23, -14, -14, -6, 9, 11, -16, 7, 20, -11, 0, -18, -23, 4, -22, -6, -11, 5, -23, 15, 3, 14, -33, 9, -34, -17, -41, -22, 29, -20, -21, 19, -1)
  );
  ----------------
  CONSTANT Layer_5_Columns    : NATURAL := 8;
  CONSTANT Layer_5_Rows       : NATURAL := 8;
  CONSTANT Layer_5_Strides    : NATURAL := 2;
  CONSTANT Layer_5_Activation : Activation_T := relu;
  CONSTANT Layer_5_Padding    : Padding_T := same;
  CONSTANT Layer_5_Values     : NATURAL := 32;
  CONSTANT Layer_5_Filter_X   : NATURAL := 3;
  CONSTANT Layer_5_Filter_Y   : NATURAL := 3;
  CONSTANT Layer_5_Filters    : NATURAL := 48;
  CONSTANT Layer_5_Inputs     : NATURAL := 289;
  CONSTANT Layer_5_Out_Offset : INTEGER := 3;
  CONSTANT Layer_5_Offset     : INTEGER := -1;
  CONSTANT Layer_5 : CNN_Weights_T(0 to Layer_5_Filters-1, 0 to Layer_5_Inputs-1) :=
  (
    (-52, 41, 10, -12, 12, -44, 14, -39, -43, 12, 15, 16, 28, 28, 4, 35, 11, -15, -8, -3, 0, -9, 0, 46, 2, 29, 21, -27, 45, 11, 11, 24, -61, 11, 6, -22, 18, -15, 65, -10, 25, -27, -6, 59, 39, 10, -42, 52, -21, 21, -1, -15, -22, 5, 44, 38, 18, -5, -18, -11, 75, -12, 23, 32, -19, 26, 20, -62, 17, -9, 29, -13, 10, -6, 1, 11, 13, -6, -48, 0, -52, 6, 15, -36, -6, -6, 12, 12, -16, -34, -8, 23, 32, -39, -20, -5, -31, 11, -6, 30, 13, 14, 15, 7, -7, 15, -53, -26, -28, 12, -15, -16, -13, -72, 59, 14, 13, -29, -24, 10, 48, -26, -13, -48, 53, -50, -22, 24, -9, -17, -41, 61, -8, -3, 29, -28, 21, 14, -53, 28, 8, 14, -55, -6, -33, -32, 1, 25, 21, -15, 42, 30, 48, 7, -17, -3, 35, -1, 16, 32, 30, 16, -17, 67, -7, 20, 10, 19, 49, -19, -51, 18, -2, 14, -79, 32, -58, 3, -5, 28, -1, -27, 0, 30, 21, 4, -36, 21, -15, 9, 11, 16, 17, -19, -19, -27, -52, 7, -37, -16, -17, -31, -62, 6, 6, -50, -22, -16, -44, -20, 31, 44, 13, -2, -20, -3, -11, -41, 11, 15, -41, -28, -60, -37, 77, 0, -18, -3, -4, -8, -30, -20, -5, -47, -52, -12, -33, -16, 32, -19, -36, -19, 65, 64, 11, -12, 8, -37, -29, -36, 6, -44, -17, -7, -28, -22, 63, 9, -25, 28, 10, -52, 0, 10, -15, -35, -7, -14, -31, -25, 38, 25, -13, -1, 12, 39, -5, 6, 13, -56, -34, -32, 36, -11, 0, -14, -35, -20, -8),
    (-21, -24, -43, 3, 21, 17, -39, -17, -12, -36, -15, -31, -24, 8, 1, 37, -36, -40, -5, -9, 17, 36, 33, -31, 17, -8, 55, -7, 20, -6, 11, 14, -5, 8, -65, 23, -5, 53, -40, -6, 8, -76, -10, -24, -8, 20, -2, 37, 0, 48, -31, -37, 8, 40, -51, -18, -6, -3, 37, -19, -4, 16, 2, -1, -4, 22, -39, 31, 2, 4, -22, 4, 7, -29, 13, 26, -21, 19, -24, 5, 38, 31, 1, -13, 2, 23, -35, -8, -14, 14, -11, -17, -22, -1, -4, -19, 33, -20, -27, -12, -21, 58, -71, -23, -51, -10, -12, -27, 0, -8, -2, 29, -13, 40, -16, -43, -10, 19, -30, -16, 21, -10, 47, -1, 43, -30, 12, -16, -5, 15, -19, -12, -27, 56, -69, -23, -47, -45, 12, -54, -30, -30, -4, 50, 19, 51, -43, -61, -11, 74, -17, -31, 16, 5, 62, -17, 13, -8, 49, -37, -28, 7, -55, -64, -2, 26, -42, -17, -1, -45, -17, -17, -21, 1, -34, 10, 9, 50, -25, 2, 0, 46, -45, 0, 13, -17, -1, -2, 6, 31, 51, -31, 2, 14, 32, -7, -5, 36, -39, -20, -40, 18, -14, 25, 28, -23, 4, -7, 10, -7, -49, -11, -17, 15, -32, -6, 38, -20, 4, 33, 11, -4, 1, -26, 3, -10, -9, -26, 4, 55, -34, -54, -76, 15, -10, -4, 24, -41, -18, 3, 15, 44, 2, -24, -12, 33, -13, -12, 29, 2, 3, 31, 1, 6, 9, -21, 17, -10, -42, -27, -30, 27, 1, -38, -34, 30, 27, -35, 7, -4, -27, 28, 32, 61, 1, 29, 26, 16, -8, 6, -1, 2, 8, -20, 18, -3, 14, 2, -2),
    (25, -44, 23, 7, -29, 8, -18, -3, -20, 3, -5, -9, 13, -11, -54, -29, -22, -7, 2, -10, 5, -45, -2, 3, 40, 52, 24, 24, 25, -14, 26, -7, 50, -51, -41, -36, -24, -15, -54, -53, -23, 8, -5, -8, 12, 16, -6, 10, -1, -8, 4, -19, 16, 1, 19, 12, 59, 26, -7, -9, 6, -37, -3, -20, -5, -30, 1, -30, 19, -51, -14, 16, -13, -3, 8, -2, 16, 30, -3, 15, -18, -13, -43, -18, 11, 19, 15, -10, -27, 39, -7, 3, 31, -24, -11, 5, 6, -56, 55, -26, 10, -3, -7, -2, -22, 9, 3, 13, 5, -4, -89, -32, -80, -11, -6, -3, 14, -28, -27, 21, 70, 39, -9, 39, -22, -68, 20, -15, 46, -73, 26, -61, 19, -13, -10, -48, -56, 28, -5, 26, 22, 0, -62, -46, -57, -2, -1, -37, 16, 0, -75, 34, 39, 9, 36, 50, 12, -57, 21, -30, 13, -35, 10, -1, 31, -36, 5, -22, -25, 16, 26, -6, 35, -9, -18, -16, -10, 17, -7, -52, 12, -6, -9, -3, -9, 35, 0, 9, -7, -32, 4, 7, -19, -23, 68, -15, -7, 9, -4, -7, -9, 19, -24, 41, -8, -27, -38, -41, -68, 5, 43, 17, 17, 0, -21, 12, -19, 25, -11, 51, -6, 8, 8, -19, -10, -28, 53, -9, -19, 11, 37, -43, 1, 30, -1, 26, -8, -29, -5, -21, -65, 12, 51, -14, -10, -28, -37, 22, 39, 31, 12, 59, -16, -17, 1, -23, -6, 0, 36, -13, 23, 23, 34, -32, -7, 8, 7, 23, -25, -21, -2, 25, -53, 24, 34, -53, -26, -12, -10, 21, 3, -14, -16, 32, 1, -12, 13, 4, -5),
    (-11, 39, 21, 46, -20, 20, -40, 39, -27, -1, -23, -24, 16, 40, -21, -12, 57, -37, 12, -15, -24, -17, 50, 20, -1, 27, 19, -46, 23, 2, -37, 9, -17, 42, 23, 34, 23, 16, -19, 36, -24, -46, 13, 26, -3, 62, -6, 9, -2, 16, -36, 24, -18, -16, 11, -8, -2, 10, -26, 46, 42, -41, 3, -18, 15, -10, 30, -21, -25, 29, 20, -8, 32, -81, -16, 97, -37, -1, 0, 0, 5, 10, -44, 8, 5, 16, 0, -7, 2, 25, -33, 53, -18, -6, 20, 10, -42, 27, 19, 44, -2, -34, 2, 29, -56, -11, 61, -29, 8, 15, -35, -31, 36, -17, 1, -32, -20, -61, 37, -2, 11, 14, -23, -28, 41, -26, -13, 45, -29, 21, 58, -24, -4, -21, 1, 40, -33, -88, -3, 13, 11, 31, 26, 21, 57, -46, 16, 10, 16, -4, 57, -22, 21, -26, -27, 11, 26, -4, -16, 23, 2, 0, 19, -47, -14, -15, 34, 45, 0, -40, -5, 12, -57, 6, -3, 6, 19, -12, 19, 20, 4, 5, 20, 18, 32, -38, -30, 2, 18, 12, 19, -20, -3, 22, -40, 28, 7, 22, 28, 1, 39, -34, 5, 29, 12, 10, -38, 7, -34, 59, -48, -27, 19, 15, 8, 38, -2, 4, -42, -31, -2, 0, -31, 43, -34, -13, -23, -11, -11, -6, 34, 7, 58, -5, -9, -2, -5, -35, -9, 8, 34, 25, -17, -38, -7, 2, 42, 29, 23, -1, -14, -29, 49, 31, 3, 44, 13, -23, -3, -21, 4, -47, 48, 11, 18, -12, -15, 13, 12, -48, 2, -27, 43, -24, -28, -81, 32, -10, 35, 25, 10, 18, 2, -3, 24, 45, 30, -50, -2),
    (-67, 10, -20, -6, 35, -22, 25, 14, -37, 19, -20, -22, 16, 10, -18, 23, 18, 16, 5, 14, -23, 19, 9, 1, 39, 35, 47, -29, 33, -4, 16, -11, -73, 11, 18, 23, 20, 15, 6, -8, -55, 35, -50, 22, 3, 22, -63, 21, 31, 34, -35, -31, 15, -5, 59, 32, 67, -6, 10, -18, 23, -19, 9, 0, 1, -37, 13, -2, -11, 13, -27, -6, -5, 0, -26, 37, 4, 37, 16, -22, 1, 22, 0, -21, -17, -34, 42, 20, 22, -15, 25, -13, 20, -38, -10, -13, -9, -28, 13, 2, -21, 34, 23, 10, -30, 1, -16, 49, 41, -15, -23, -32, 18, -4, 7, -18, 30, 8, -29, 47, 20, -5, -27, 22, -2, -1, 37, -30, 10, -44, 9, 12, -18, 3, -22, -59, -17, 27, 12, 3, 6, -35, 20, -44, -56, -2, 20, 51, -11, -9, -12, -25, 20, -21, 15, 26, 5, -25, -6, 21, 5, 3, -6, -19, 0, -14, -38, -12, 26, -30, -2, 5, -20, -1, 1, -11, -17, 14, -26, 61, 48, -1, 1, -1, -21, 11, 12, -26, 20, -35, -40, 1, -5, 18, -3, -23, 19, -34, -45, -16, -20, 26, -6, -3, -24, -41, -24, -21, 11, 6, 42, 0, -3, -46, 22, 16, -6, 3, -36, 2, -12, -33, -10, -53, -4, -11, 10, 32, 18, -42, -50, 1, -38, 18, 11, -52, -49, 29, 57, 35, -47, 2, -5, 31, -21, -6, 45, 20, -38, -60, 30, -26, 64, -15, -29, -32, -16, -17, 9, 7, 43, 41, -24, -6, 0, 0, 18, -44, -41, 35, 53, 9, 16, -5, -1, -31, 14, 44, -22, 27, 11, 31, 43, -28, 39, 2, 22, -9, -5),
    (19, -28, 31, 41, 21, 22, -2, -26, -23, -13, -25, -29, -42, 26, 44, -8, -31, -79, -6, -66, -30, 15, 67, 44, 2, 7, -7, 13, 37, -44, -49, 41, -16, 7, 12, 28, 28, 14, -10, 3, -30, -49, 2, -19, -5, 42, 31, 8, 8, 9, -45, -64, -33, 41, 29, 43, -28, -14, 17, -9, 37, -10, -48, 18, -26, 13, 19, 20, 3, -4, 5, 34, 3, -54, 25, 16, -17, 42, 28, 18, 4, 1, -55, -43, -22, 42, 14, 33, -30, 23, 7, -39, 19, -9, -42, 10, 52, -25, 22, 57, -59, -32, 59, 9, 33, -6, 31, 14, -14, -5, -18, 3, 8, -52, 15, 9, 8, -4, 39, -11, 45, -39, -26, -2, 24, 32, 10, -1, 32, -30, 34, 8, -11, -8, 52, 29, -19, -7, 21, -45, -42, 37, 31, -12, 4, -19, 27, -11, -36, -7, -32, -15, 9, -11, 1, -31, 38, -4, 4, 47, 9, 5, 22, 11, -15, 24, 18, -6, -39, -58, 9, -29, -20, 11, 18, 25, 20, -16, 14, 4, -14, 35, 19, -35, 16, 6, -2, -29, 34, 10, -14, 22, -12, -16, 9, -16, 11, -34, 39, -24, 24, 30, -10, 35, 29, -47, -58, 1, -23, 24, -20, 26, -20, -3, 52, 28, -15, -43, 7, -6, -15, 41, 20, -29, 40, -43, -17, 12, 11, -2, 55, -38, 7, 42, 4, 41, 34, -54, -52, -2, -16, -3, -34, 20, -8, 31, 37, 53, 11, -25, -20, -6, 43, 48, 18, 37, 28, -11, 23, -13, -42, -34, 30, -15, -30, 47, -62, 4, -34, -26, -23, -27, 1, -22, -14, -2, -14, -4, 48, -21, 19, -32, -10, -44, 11, 18, -16, 23, 16),
    (-8, 4, -16, 8, -13, -9, -59, -3, 8, -17, -5, 38, -25, -16, -79, -14, 28, 10, -23, 14, 12, -50, 4, 12, 2, 16, -24, 22, -8, 1, 30, -16, 12, -27, -35, 14, 35, -26, -46, -17, 3, -20, -12, 6, 21, 34, -87, -23, -31, -15, -45, -39, 14, -16, 26, 25, 11, -4, 18, -7, 32, -34, -18, 13, 16, -19, -16, -7, 25, -4, 9, -26, 11, -34, -28, 10, 32, -10, -63, -20, 49, 24, -22, -33, -1, -20, -23, 7, 23, 4, 26, -19, 5, -2, 37, -29, -7, 26, 24, -21, -34, 40, 12, -28, 21, 2, 2, 0, -17, -3, -22, 17, 18, 25, -57, -7, 32, -2, 53, -11, 37, -23, 20, 11, 65, 9, 13, -4, 61, -37, 25, -11, -8, 33, 0, -66, 12, -7, -45, 25, -4, -40, -25, 43, -52, 46, -58, -13, 17, 11, 2, -14, 50, -37, 3, 29, 27, 25, 48, -16, 8, -5, -58, -13, -18, 26, 7, -52, -18, -5, -43, -1, -32, -40, -18, 43, -19, 13, 1, -6, 27, 11, -17, 23, 26, 11, -3, 30, 3, 24, 15, -30, 13, 15, -48, -40, -6, 58, -23, -26, 11, -5, 22, 10, 6, 11, 22, 14, -23, 13, -23, 34, 15, 59, -2, -32, 22, -28, 23, 5, 15, -8, 2, -56, 51, -15, 3, -28, -2, 67, 2, -37, 24, -6, -17, 6, -15, -3, 24, 25, -13, 51, -26, 11, 15, 43, -59, -28, 21, -25, 19, 30, -7, -4, 9, -34, 54, 21, 6, -22, -48, 28, -16, 1, -25, -2, -40, 7, -12, 12, 17, 1, 23, 50, 25, -8, 7, 26, -54, 6, 9, 8, -17, 2, -41, -24, -12, -11, -3),
    (-9, 11, 29, -29, -47, -6, 1, 34, -20, -49, 11, 47, -42, -4, 27, -23, 26, 28, 7, -49, 11, 12, 20, 3, -7, 13, -5, -61, -4, -37, 1, -28, -4, -20, 44, 25, 4, -39, 28, 7, -18, -34, 3, 12, -34, -9, -57, -25, 42, 4, -28, -17, 15, -25, 16, -14, -24, -24, -27, 5, 50, 27, 21, 9, -28, -69, 28, 26, -14, -9, 20, -37, -43, -3, -49, -30, 2, -11, -42, -1, -1, 6, -2, -45, -19, -1, 8, -57, 11, 3, -22, -7, 3, 54, -10, -40, 4, 25, -44, 18, -10, 45, 13, 13, 55, -16, 18, 1, -18, -23, -40, 7, 25, 28, -41, -7, 31, 39, -27, 7, 22, 3, 4, -8, 60, 36, 34, 12, -10, 18, -26, -10, -38, 17, 37, -55, 43, -8, -12, 33, -13, -27, -67, 50, -3, 12, -44, 6, -13, 9, 20, 59, 16, -29, -9, -4, 58, 46, 54, -44, 28, -32, 20, -2, -26, -13, 69, -15, 49, -26, 46, 49, -12, 16, -12, 8, -21, 20, 8, 45, -20, 9, -3, 11, 33, 20, 1, -1, 71, 41, -7, 2, 30, 15, -13, -6, -12, 3, 7, 10, -21, 20, -17, -18, -38, 11, -50, 16, 0, 4, 6, 14, 6, -5, -23, 29, -34, -46, 14, 21, 7, -2, -25, 24, 31, 2, 5, 4, 2, -11, -27, -41, 29, 29, -20, -7, 8, -8, -53, 8, -40, 22, 16, 26, 2, 2, -10, 19, 34, -24, 32, -5, -28, 1, -2, -17, 28, -28, 5, -25, 4, -1, -43, -5, -15, 11, -45, 13, -9, 6, -46, 27, -6, 0, 16, -10, 24, 26, -17, 26, 25, -14, -7, -9, -21, 19, 5, -16, 3),
    (-12, -29, 9, -16, 6, 16, -23, -34, -3, -34, -34, 31, -20, 36, -13, 2, -8, -11, 48, -7, 21, 42, -9, -14, -5, 22, -2, 32, -57, -42, -39, -4, -12, -3, -15, 5, -9, -46, -25, -4, 17, -49, -60, 60, -40, 12, -38, 0, -10, 1, 54, 0, -10, 30, -16, 4, -21, 20, 0, 36, -77, -45, -24, 61, 12, 3, -9, -5, 14, -28, -51, 6, 4, -28, -47, 39, -57, -26, -13, -26, 11, -4, 15, 15, -6, 20, -22, 0, -8, 10, -2, 2, -38, -11, -22, 23, -23, 10, 6, 42, -1, 23, 2, 7, -60, -14, 18, -6, 21, 34, 38, 25, -9, -5, -24, -21, -14, 29, 36, 33, -20, 7, -2, -1, 64, -51, -55, 44, -35, 35, -7, 45, 11, -6, 20, 36, -45, -26, 2, -24, 10, 31, 45, 38, 20, 14, -34, -66, -8, 17, 23, 55, 9, 10, 16, -21, 72, -5, -19, 44, -16, 30, -3, 19, -11, -22, 45, -7, -43, -19, -10, -26, 35, 44, -19, 66, 29, 29, -44, -54, -17, 8, -2, 43, 13, -3, 1, 25, 74, -14, 14, 27, 42, -41, -21, 28, -51, 17, -6, -20, -9, -3, -10, 3, -1, -5, 1, -44, -35, 3, 28, -13, 41, 7, 11, -18, 15, -20, -7, -21, 19, -7, -10, 6, 42, -18, -42, 41, -11, 14, -7, -13, 34, -4, -27, -25, -1, -23, -42, -26, -8, -53, 30, 26, 31, -5, 12, -17, 41, -9, -16, -6, 29, 23, 4, -5, 25, -7, -9, 13, -6, -43, -31, -20, 40, 11, -21, -14, 7, -54, -40, -27, -28, -13, -4, 36, -11, -53, 5, -26, 27, -12, -21, 1, -26, -4, 9, -36, -3),
    (33, 34, -16, 27, -34, 17, 56, -10, -6, 31, 49, -28, 12, 3, 10, -41, -57, 19, -38, -32, -8, -6, -28, -41, 20, -48, 18, -26, 34, 36, 5, -17, 2, -33, -20, 14, 22, 4, -12, 22, 29, 25, 23, -33, -1, 8, 60, 3, -25, 23, 30, -22, -1, 29, -30, -20, 17, -20, 1, -37, 9, 53, -19, 30, -15, 24, 14, -31, -39, -13, 21, -25, 5, 10, 5, 23, 24, -3, -23, 47, 42, 15, -21, 18, -28, 21, 0, 14, 11, -2, -24, -28, 28, 30, 2, -6, -33, 17, -38, 43, 9, 24, 18, 20, 1, -45, 53, -10, -29, 11, 22, -3, 17, -27, -28, -19, -8, 17, 3, -1, 3, -4, 12, 12, -7, 39, 8, 35, -3, 61, -2, 11, -42, 64, 52, -10, -19, -13, 58, 0, -19, 3, -52, 1, 51, 31, 9, -27, -24, -5, 30, -9, 4, -10, 4, 9, -3, 44, 0, 54, 27, -11, 11, -61, -5, -48, 11, -7, -9, 29, -46, 24, -11, 8, 28, -30, 21, 29, -20, 33, -4, -16, 74, -65, -37, -14, -47, 41, 44, -5, 11, -31, 16, -20, -19, -13, 34, -20, 36, -11, 25, 4, 18, 7, -40, -40, -101, -14, -9, 37, 19, -19, -21, 30, -27, -11, -47, 3, -40, 74, -39, 23, 26, -19, -1, 21, 27, -8, 1, -57, 30, -19, -8, 18, 30, -20, 11, -113, -40, -40, 47, 35, -33, 2, -23, 3, 36, -19, 13, -22, -20, 54, -5, 24, 20, -3, 29, -35, -17, -66, 7, -23, -23, 26, 37, 29, 34, 8, 13, 4, -1, 26, -6, 7, 5, 43, -13, -43, 5, -18, 13, 8, -48, -29, -50, -11, -51, -68, 13),
    (-16, 49, 18, -12, -28, -3, 6, 21, -12, -30, 1, -27, -31, -11, 25, -1, 17, -41, -6, 14, -5, 29, -27, -30, 7, 16, -8, 6, -19, 9, 17, -8, -14, 32, 32, -20, 23, 6, -22, 2, -26, -32, -3, 14, 6, 13, 37, -23, 40, 64, 1, 11, -35, -9, -9, -16, -9, 24, -22, 10, -17, 0, 14, -21, -31, 31, 9, 1, 0, -31, -68, -21, -40, -25, 9, 33, 7, 2, -7, -7, 4, 72, 0, -2, -18, 20, -42, -4, 1, 12, -10, 42, 2, 13, -12, -51, -25, 45, -8, -1, 8, 21, -17, 31, -21, 11, 35, 9, -15, -10, 24, 19, 54, 6, -13, -59, 17, 33, -2, -29, -2, 3, -23, 11, -19, -7, 18, 42, -44, 73, 2, -67, 10, 36, -21, 53, -39, -38, 48, 20, -19, -14, 40, 21, 92, 67, -19, 11, -1, 24, -30, -73, -7, 43, -41, 18, 10, 4, 46, -24, -18, 54, 25, -38, -16, 9, -73, 16, -44, -27, 27, 30, 17, -6, 16, -22, 34, 61, -18, 36, -18, 8, -28, -11, 27, 41, -18, 43, 34, -18, 3, -75, -43, 6, 28, -3, -13, 19, -22, 7, -10, 14, 25, 8, 0, -18, 4, -6, -5, 34, 14, -78, -6, 13, 42, 16, 8, -11, 14, -5, 10, 11, 9, -18, -57, 38, 0, 2, 9, 20, -24, 13, 19, 14, 23, 2, -8, -23, -49, -5, 43, 21, -26, -41, 26, 38, -22, -22, 2, -5, 8, -20, 34, 40, 46, 18, -8, 56, -7, -61, -35, -15, -4, -6, -16, 11, -8, 18, 29, -21, -5, 7, 43, -9, 4, 4, -25, -5, -4, -35, 18, 13, -33, 3, 38, -20, 8, -49, -12),
    (13, 3, 7, 30, 16, -7, -19, -26, 1, 15, 18, 54, 2, -49, -44, -30, -12, 30, 25, 29, 13, -15, -63, -24, 17, -15, 0, 46, -41, -47, 24, 17, 61, -48, 29, -17, 43, -6, -12, -32, -3, 66, 2, 35, 33, -40, -10, -14, -62, -10, 29, 58, 36, 12, -25, 3, -17, -4, -27, 40, -53, 1, 22, 0, 36, -15, 15, 2, -2, -15, -30, -42, 14, 21, 14, 12, 20, 24, 31, -31, -50, -8, -8, 39, 56, 31, -16, 39, -5, -18, -22, -11, 12, 28, 3, 6, -8, 30, 15, 11, -37, -18, 37, -29, 35, -11, 57, 29, -26, -27, -8, -37, -26, 26, 16, 45, 23, -7, -45, -29, -1, 6, -27, -1, -27, 37, 24, -31, 60, -4, 20, -45, -17, 7, -20, -58, 4, 60, -4, 11, 48, -45, -32, -18, -35, -29, 4, 65, 47, -19, -2, -18, 4, -22, -48, 30, -58, -32, 23, -57, 49, -23, -8, -32, 13, 46, -23, -1, 1, 34, -19, 0, 23, -5, 25, -8, -18, -12, -25, 51, 59, 35, 17, 10, 2, -36, -37, 13, -18, 18, 5, -41, -7, 67, -16, -9, -9, -2, 15, 27, 51, -12, -4, 4, -17, 18, -5, 6, 19, -2, -1, -27, -7, -14, 8, -21, -38, -32, -8, 27, -14, 27, -14, 5, 2, -1, -17, -30, -16, 20, -39, -20, 44, -1, -8, 37, -5, -23, -34, -18, 21, 32, -18, 0, 14, -24, 4, -20, 25, -10, -24, 32, 6, -10, 4, -31, 15, 9, 2, -38, -5, 1, -55, -21, 9, 33, -22, 17, -5, -11, 15, 26, 27, -27, -18, 26, 10, 31, -5, -8, 12, 0, -16, 15, -14, -21, -9, -50, -19),
    (7, 41, -42, -11, 2, 6, 2, -16, 26, -46, -18, 14, -5, -41, -26, 21, -1, 36, 7, 48, -50, -25, 40, -25, -14, 34, -3, 51, -21, -14, -42, -40, -15, 20, -8, -28, -10, -3, -27, -36, 6, 50, -26, 38, 45, -19, 2, 21, 4, 36, 19, -33, -23, -9, -14, 31, -31, 3, -15, 89, -29, -4, -25, -6, -3, -36, -8, 32, 29, -27, 9, 26, -23, 54, 3, 6, -4, -31, 15, -35, 6, 0, 16, -48, -3, -37, 18, 49, 35, -10, -8, -13, -21, -13, -16, 12, -13, 66, 4, -54, -24, -5, 4, 37, 1, 4, 49, 52, 13, 0, -1, 44, 16, -31, -19, 22, -20, 34, 26, 30, -49, 9, -30, 5, -18, -56, -30, -16, -42, 61, 37, -7, -4, -22, 7, -7, -24, 71, -12, 78, 27, 1, -28, 32, -1, 15, 6, -27, -6, 21, -48, 51, -12, 51, -12, 83, -31, -8, -15, -15, -52, 3, -11, 7, 17, -45, -44, -5, -91, 12, -38, 10, 24, -23, 0, -30, -18, 12, 28, -54, -40, -6, -26, 5, 19, 8, -21, 34, -3, 11, -12, 6, -16, 29, 24, -13, -33, -2, 20, 30, 15, -28, 30, 55, 16, -2, 17, 30, 9, -10, 21, 14, 20, -38, -13, -10, 1, -26, 12, 16, -19, 17, 6, -12, -22, 27, 38, 14, -9, -38, -6, 28, -26, 29, -7, 27, 14, -26, -31, 12, -2, 32, 28, -12, -8, -31, -26, 38, 16, 31, 3, 34, -18, -22, 11, -8, 9, 3, -30, -11, -26, -11, -71, -17, -20, -7, 23, -31, -1, 30, 19, 10, -6, 18, 43, 48, 7, -27, -42, 0, -30, 4, -37, 36, -12, -41, -15, -1, -8),
    (-31, 42, -1, 18, 6, -14, -11, 46, 7, 1, 39, -50, -11, 6, 46, -20, 32, -41, 40, 15, -33, -40, -13, 6, -29, 9, 28, -6, -52, -21, -27, 5, -41, 51, -9, 11, 0, -64, -14, 38, 24, -39, -3, -56, -25, -9, 56, 22, 18, -27, 44, -17, -26, -7, -21, -20, -25, -15, 20, -27, -25, -52, -59, 27, -6, 38, 25, -3, -6, -56, -21, 46, 12, -28, 9, -44, -36, -11, 42, -19, 3, 14, 31, 11, -20, 2, -43, -26, -4, -30, -3, -43, -45, -12, -44, 12, -67, 19, 42, -9, 40, 15, -23, 8, -50, -16, 7, -22, 16, 33, 26, 20, 22, -17, 22, -48, -14, -5, -3, 12, 33, 39, -10, -19, 53, 39, 15, 8, -102, 3, 47, 22, 31, -33, -2, 34, -20, -45, 36, -3, 14, 19, 10, 44, 63, 9, -4, -81, 12, -16, -3, -2, 39, 17, -20, -44, 53, 20, -11, 60, -90, 17, 34, 49, 24, -31, -23, 32, -28, -28, 27, -34, 1, 21, -5, -4, 79, 35, -6, -58, -24, -9, -41, 40, 22, 19, -10, -41, 8, -18, -2, 39, -16, 12, -10, 56, -22, -22, 6, -9, -32, 6, -1, -1, 12, -18, 0, -16, 0, 47, 5, 32, -4, 10, 9, 2, 6, -23, 16, 7, 81, 2, -10, 23, -19, -35, -19, 72, 19, 13, -7, -6, -31, -7, 45, -19, -9, -13, 11, -2, -61, 31, 8, -9, -3, 19, -36, -16, 15, 25, 18, -16, 55, -28, -6, 30, -20, 4, 33, 59, 8, 4, -31, -24, 0, -2, 29, 15, 6, -14, -33, 23, -9, 29, -20, -5, -16, 24, -35, -7, -5, 38, -43, -1, 21, -25, 35, 58, -7),
    (-12, -20, 34, 10, -10, -26, 27, 18, 12, -27, 19, -3, -40, -51, -20, -31, -25, -69, 19, -20, 19, -11, 31, -30, -14, -26, -21, 20, 18, 5, 31, 25, 41, -13, 29, 21, 5, -23, -9, -29, -3, -19, -17, -1, 25, -25, -1, -42, -59, -14, 37, -10, -40, -6, -17, -6, -29, -24, 22, 12, 13, -19, 15, 46, 6, 5, 5, 20, 40, 9, -52, -25, -15, -12, -14, 7, 24, -13, 2, 24, -16, 18, 41, -7, -15, 10, 11, 2, -11, -13, -16, 16, -10, 38, -38, 17, 11, -49, 34, 21, -24, -37, 32, -17, 58, -1, 4, 16, 17, -51, -76, 14, 19, 10, -94, 18, -25, 16, 65, 59, -24, -13, -1, -39, -5, 28, 24, 25, 15, -44, 45, 7, -3, -38, 71, -16, 51, 15, 17, 34, 3, -46, -69, -26, -8, -32, -41, 41, -6, 2, 43, 48, 50, -9, -13, -27, 53, 54, 40, 32, -16, -21, 20, 7, -33, -41, 15, -4, -15, -7, -1, -9, -17, -26, 0, -25, 6, -15, 24, -5, -24, 4, 7, 49, 23, -50, -26, 19, 32, -6, 11, 3, 8, 1, -10, -9, 28, -7, -63, -20, -12, 13, -6, -4, -2, 13, 26, 3, -16, 43, 13, 4, -21, -21, 10, 8, 0, 9, 7, 3, 12, -36, -8, 21, 45, -59, 15, 26, -5, -23, -8, -31, 25, 83, -26, 43, 11, -26, -16, 12, -50, 26, -28, 37, 14, -16, 15, 42, -18, -11, 6, -14, 20, 31, 38, -35, 44, -66, -2, -1, -2, -13, 45, -21, 8, 64, -19, 14, -1, -48, -29, -6, -18, 14, -38, 7, 28, 7, 5, 49, 12, -30, -44, -10, -2, 24, -23, -8, 12),
    (-23, 9, -20, -30, -21, 15, 45, -2, 39, -40, 7, 16, -1, -17, 11, -23, 27, 42, 57, -51, 2, -43, -65, -19, 39, 15, -21, 60, -15, -3, 23, -2, -47, -26, -1, 18, 3, -5, 67, -5, 2, -12, 42, 20, -6, -9, 3, -16, -18, 3, 43, 7, 24, -36, -35, 4, 27, 5, -11, 70, -26, -34, 4, -6, 5, -13, -27, 16, 25, -21, 45, -4, -29, 2, 21, -6, -2, -6, 22, -34, -5, -13, 15, -5, 13, -35, -6, -13, 3, 15, 17, 5, -19, -27, 11, 29, 16, 55, -8, 34, 7, -27, 53, 3, 54, -33, 38, 60, -7, -14, 0, 10, 25, 33, 58, 8, 11, -13, -75, -27, -21, 7, -17, 63, -62, 2, 7, 31, 18, -11, -33, 51, 13, -9, 85, 3, 49, -2, 39, 57, 8, -10, 10, -50, -63, -31, 74, 28, 7, -76, -96, -4, -17, -26, -31, 63, -75, -12, 11, 41, 22, -25, -13, 52, -8, -14, 46, -10, 11, -1, 35, 25, 4, -11, 0, -33, -37, -31, -5, 23, 15, -31, -21, 0, -6, -5, 6, 35, -29, -6, -13, 17, 15, 1, 2, 23, 0, -19, 24, 11, 42, -31, 27, 7, -15, -11, -30, -13, 30, 31, 44, 19, -4, -20, -43, -11, -21, -34, 2, -15, -18, -6, 1, 37, 62, 4, 12, 35, -15, -13, 12, -11, 15, 4, 14, 35, 28, 3, 10, -51, -2, -8, 42, 34, 14, -43, -84, -11, -37, -3, -2, 31, -71, 9, 0, 19, 17, -12, 15, 0, 7, 15, 9, -6, 21, 5, -9, 3, 14, -13, -4, -12, -21, 11, 7, 32, 11, -19, -29, -5, -9, 15, -18, 34, -33, 0, -13, -18, -9),
    (21, -31, -2, 59, 20, -16, 0, -8, 11, -26, 37, 7, 15, 8, -26, -5, -86, -45, 18, 44, 18, 12, -59, 10, -18, -6, 23, 13, -45, -7, -15, 19, -4, -50, -25, 34, 3, 2, -20, -2, -12, -25, 52, -73, 8, 24, 26, -37, -16, -31, 30, 13, -13, 64, -10, 2, -20, -4, 12, 9, -67, -52, -37, 67, -5, -22, -45, -56, -4, -42, 25, 7, 17, -28, 82, -72, -67, 11, 16, 1, 1, 22, 16, -64, -34, 28, -24, -19, 4, -8, 19, -67, -9, -27, -51, 1, 72, -70, 8, 25, 8, -15, -8, 26, 7, -26, 27, -73, -2, 16, -1, 6, -76, 15, -9, 10, 20, 22, -15, 1, -41, 26, -4, 31, -64, 8, -45, 69, 11, 9, -22, 44, -15, -27, -5, 37, -23, -36, 48, -17, -5, 37, 17, 21, -28, -47, -3, -90, 1, 51, 3, -6, 15, -12, 0, -22, 3, -35, -47, 95, -63, 21, -9, -33, -12, 47, -2, 58, -4, -39, 48, -36, -40, 27, 0, 14, 49, 43, 10, -42, -26, -20, 24, -41, -7, -32, -3, -73, 29, -31, -1, -2, 33, -8, 13, 7, -27, -2, 19, -12, 40, -2, 43, -27, 15, 10, -4, 4, 13, 10, 3, -58, -11, -4, -54, 20, -24, -24, 2, -9, 33, -7, -23, 49, 1, 28, -55, 25, 3, 11, 41, 49, 50, -53, 41, -27, 21, 18, 2, -15, 1, -5, -15, -94, -21, 0, 7, -1, 3, -18, -25, -9, 15, -4, -5, 35, -52, 3, -38, 8, 26, 5, 17, -40, 3, -27, -7, -3, 9, -16, -17, -10, 16, -19, -14, -12, 3, -21, -51, 0, 61, -5, -9, 31, 14, 3, 23, 12, -4),
    (6, -22, 11, 24, -20, -16, 53, -8, -17, 50, -33, 28, 20, -45, 0, -15, -12, -57, 28, 2, -9, -21, 16, 10, 3, 23, -15, 27, -52, -18, 23, 24, 35, -11, 13, 35, -16, 14, 25, -80, -31, 19, 13, 24, 56, -24, 4, 2, -22, -16, 33, -23, 1, -9, -54, 14, 22, 10, 5, 18, -34, -11, 22, -11, 13, -27, 0, 10, -1, 13, -17, -32, -18, 18, 14, 20, 56, -30, 12, 26, -37, 11, 23, -18, 6, 21, -13, 21, 29, 18, -1, 26, -39, -11, -30, 11, -2, -15, 54, 23, -19, 20, 70, 22, -43, 28, -7, 20, -1, -70, -40, -36, -30, -22, 49, 1, -11, -45, 8, 0, 39, 40, -16, 29, -38, 27, 10, 10, 43, -33, 46, 7, -4, 19, 65, -44, -45, 62, 58, 32, 31, -73, -67, -1, -32, -15, 11, -13, 30, -36, -19, 12, 70, 27, -26, 44, -29, -7, 24, 21, 25, -43, 0, 23, -24, -16, 20, -75, -28, 29, 0, 46, 58, -50, -46, 14, -40, -22, 12, -28, 49, -12, 3, 30, 49, 3, 5, 39, -17, -26, 3, 21, -9, -24, 4, 13, -37, -47, 37, 15, 25, -23, -3, 3, -5, -29, -31, -35, -15, -20, 19, -10, -4, 9, 2, -13, -33, -12, -38, -8, 17, 6, 3, 38, 13, -2, 36, 1, 3, -17, -3, 6, 6, 1, 4, 26, -31, -58, -79, -9, -45, -4, 15, 33, 4, -10, 42, -9, -33, 3, -52, 30, -20, -6, 29, -11, -4, -13, 1, 11, -20, 15, -14, 4, -6, 21, -20, 11, -20, -10, -41, -21, -55, -1, -3, -7, 18, -28, 43, 22, 19, 37, -6, 28, -16, -17, -12, -16, -9),
    (-36, 18, -41, -46, 31, -12, 24, 17, -18, 0, 10, -7, -1, 13, 1, 27, 12, -20, 52, -11, -21, -27, -58, -3, 28, 46, -2, 32, -26, -30, 24, -21, -47, 23, -1, -24, 29, -42, 9, 11, -44, 5, 31, -23, -28, 35, 24, -10, -5, 5, 63, -15, -25, -51, -57, -55, 42, 48, 24, 63, -43, -44, -9, -2, -45, 4, 48, -76, -35, -10, -20, -1, -2, 4, -21, -19, -43, 16, 30, -7, -16, 33, 42, 21, 0, 2, 31, -35, 22, -11, -38, 35, -10, -28, -22, -4, -20, 24, -47, -12, -8, -22, 0, -8, -31, -36, -17, 29, 28, -1, 4, 37, 24, -12, -3, -19, 27, 3, -35, -2, 39, 76, 14, 59, 1, -33, -14, 12, -94, 14, -29, 22, 3, -19, -5, -8, -62, -70, 14, -41, -7, 34, 35, 15, 20, -34, 56, -58, -41, -9, -55, -34, 50, 74, 31, 58, -18, -88, -43, 44, -73, 8, 9, -5, -23, -11, -7, 33, -54, -38, 35, -60, -38, 24, 21, 22, 13, -10, 36, 4, -14, 6, -31, -54, 23, 28, 0, 10, -28, -66, -33, 32, 2, -1, -16, -14, -3, 4, 10, 7, -44, 21, -31, 38, 14, -10, -5, -25, -9, -7, -23, -39, -5, -6, 34, 10, 33, 38, 21, 42, 13, 8, -1, 10, -39, -2, -15, 37, 24, -3, 15, 9, -67, 0, 21, 7, 27, 16, -7, 12, -8, -4, -11, -49, -11, -10, 7, -9, 25, 59, 16, 16, 22, -29, -3, 21, -24, 19, -10, 5, 15, -6, 3, 13, -30, -20, 20, 2, 22, 17, -11, 21, 17, -23, -9, -29, -2, 10, -17, -39, 11, -5, 42, 3, 35, -22, -17, 37, -7),
    (8, -13, 28, 18, -8, 9, 24, -39, -3, 73, -3, 13, 14, -22, -95, -4, -1, -6, 14, 27, 31, -3, -6, 30, 30, 37, -13, 14, 43, 20, 27, -15, 10, -8, 13, 13, -2, 24, 22, -9, 29, 25, 22, 24, 35, 32, -46, -5, -7, 3, 41, 57, 16, -13, -7, 9, 16, -26, -16, 10, 68, 9, 49, 6, 14, -14, -20, 37, -25, 15, -2, 1, 29, -15, 1, 23, -1, 9, -3, 24, -44, 10, -13, 15, -30, 1, 9, 7, 2, 7, 10, 21, 39, -17, 6, 3, 65, -69, 29, 13, 5, 0, 5, -59, 50, 72, -71, 39, 17, -43, -36, -47, -83, -32, 66, 84, 25, -37, 8, 9, 32, -5, -38, 4, -37, -26, -15, 3, 73, -27, 21, 25, -18, 8, 7, -58, 88, 29, -19, 13, -27, -10, -23, -27, -93, -37, 38, 100, 10, -4, 12, 4, -22, -16, -15, -7, 7, -16, -15, -3, 35, -18, -1, 25, -12, 9, -4, -26, 18, -6, -12, -4, -44, -5, 17, -13, -29, -18, 16, 67, -25, 14, -9, -1, -11, -36, 18, 18, 35, -11, 5, 6, 22, 11, 7, 9, -55, 26, -8, 25, -9, -12, 18, -6, 8, 22, 35, -10, -21, -19, 3, -31, -10, -25, 82, -13, -3, -3, 23, 8, -22, -46, -27, 11, 34, 6, 31, -25, 4, 20, -41, 20, -5, -46, 13, -33, 4, 17, 0, 10, -11, -25, -24, -51, -12, -9, -23, -29, -22, -39, 10, -31, -3, 5, -5, 2, 26, -31, 5, -41, -23, 5, 2, -15, -20, -17, -30, -52, -3, -20, -7, 1, 30, -1, -2, -30, -1, 1, 0, -13, -14, 16, 12, -33, 9, 40, -8, -38, -1),
    (-51, -20, -1, 22, -15, 59, 24, -5, -7, -29, 31, -2, -44, -5, 26, 16, -28, 84, 0, -1, 14, -5, -32, -10, 20, -17, -10, 21, -8, 40, 16, 2, 25, -7, -12, -23, -2, 49, -16, -45, -11, -54, 38, 28, 0, -51, 39, 15, -28, 72, -11, -15, -15, 28, -73, -50, 68, -24, 43, 41, 16, 13, 44, -30, 6, 2, -14, -30, -35, 38, -34, -12, 7, -43, -16, -22, -1, -21, 10, 19, 14, -12, 14, -4, -9, 27, -6, -26, 64, -8, -1, 22, -15, -3, -16, -44, 38, 17, -49, 14, -14, 41, -50, -26, 14, -53, -13, -33, 3, 21, -1, 1, -26, 7, -13, 6, -7, 38, -21, -10, 27, -28, 49, 13, 5, 13, 35, 0, 37, 29, -62, -40, -42, 100, -106, -33, 13, -68, -30, -17, -4, -20, -4, 8, 2, 43, 10, -13, -1, 61, -74, -64, 41, -14, 69, 18, -15, -1, 50, -20, 34, 18, 25, -16, -57, 36, -45, -21, -30, -4, 27, -13, -10, 18, -11, -8, -12, 46, -21, -9, -1, 33, -68, -28, 40, -15, 48, 44, -29, -41, 5, -23, 50, -17, -36, -59, -4, 26, -3, -18, -10, 11, 2, -10, -31, 19, -5, 2, -21, 5, -6, -35, -1, 21, 18, 0, -7, 35, 11, 1, -28, 3, -44, -21, 19, -6, -19, -46, -6, 24, 5, -10, -48, 39, -38, 10, -6, -18, -15, -20, 56, 9, -13, -71, 5, 29, -38, -3, 30, 8, 13, 15, -14, -48, -20, 7, -10, -19, 15, -37, -12, 3, -5, -7, -40, 49, 11, 43, 29, -50, -43, -24, 30, -2, -35, 2, 36, 13, 38, 16, 25, 18, -2, 29, 25, 10, 14, -78, -17),
    (-3, -7, -2, -14, -7, -26, 8, 45, 15, -41, -11, 29, -10, 1, 7, 21, 13, 3, -30, -54, -41, -7, 21, 26, -5, -6, -15, 23, 60, 7, -21, -4, 7, -54, 34, -24, 28, 20, -50, 18, -51, 43, -1, 2, -2, 9, 11, 15, 25, 69, -9, -23, 6, 25, -22, 30, 12, -2, 6, 64, 48, 8, 14, -17, -32, -2, 54, -57, 16, -13, -17, -7, -9, 13, -2, -17, -20, 34, 13, -9, 16, 6, -18, -42, 2, 23, -13, -2, 15, 3, 5, 25, 36, -13, -3, 8, -22, 51, 7, -82, -9, 24, 2, -8, 3, 5, -45, 13, 3, -10, -22, 35, 42, -46, 0, 6, 0, 0, -46, -32, 23, 26, -5, 40, -2, -34, 21, -42, 16, 0, -36, -84, -17, 45, -8, -49, -55, 43, -39, 20, -5, -28, -26, 15, 15, 69, 3, -35, -30, -43, 0, -18, 80, 18, -8, 62, 24, -29, 54, -27, 8, -46, 31, 1, -5, 55, -34, -22, -11, 53, -33, 14, -17, -13, -34, 4, 2, 43, -10, -20, 1, -1, -54, -15, 74, -11, 26, 23, 66, -53, 13, 14, -34, 5, 14, -33, -26, 28, 37, 22, -25, -18, 4, 7, 1, 6, -5, 21, 32, -26, -36, 16, 2, -2, -24, -6, 48, 19, -10, 42, 26, -13, 32, 20, 13, -4, -1, -61, -41, 12, -24, -39, -1, 11, -14, 20, -10, -13, -17, 27, 1, 15, -14, 12, 30, 11, -37, -28, 14, -3, 33, 56, -2, -41, 18, -19, 19, -13, -16, -38, -5, 30, -19, -25, -20, 7, 2, -2, -8, -44, -27, 12, -24, 32, 6, 0, 19, 7, -26, -42, 23, -34, -10, 8, -34, -52, 12, -55, -12),
    (-41, -27, -7, 6, -30, -7, -26, -1, 23, 10, 8, 13, -7, 8, -2, -25, -3, 6, 7, 22, 1, -33, -6, 43, -21, 4, -34, 0, -9, -51, -24, 32, -12, 23, -9, 13, 19, 26, -12, -17, -31, 5, -6, 16, 47, -13, -67, -32, -20, 23, 14, -12, -19, 9, -10, 20, 23, -4, 27, -4, -21, 20, 2, 21, -25, 52, 0, -2, 39, -2, -18, -20, -2, 2, 0, -11, 23, -21, -39, 13, 43, 15, -19, -1, -29, 4, 14, 14, 24, -23, -36, 17, -16, 18, -20, 0, -22, 31, 2, -2, -12, 35, -55, -3, -45, -14, -17, 19, 25, 23, 35, 36, -26, -4, 17, -41, -2, 39, 37, 11, -26, 9, -5, -4, -5, -4, -3, -2, -104, 85, 0, -19, 11, 18, -22, 33, -80, -57, -27, 24, 29, -20, 13, 20, 62, 32, 0, -79, -32, 36, -35, 28, 25, 6, -30, 7, 10, -8, 13, 35, -53, 44, 56, -13, 5, -39, -19, 23, -21, 2, 32, 0, 24, -40, -9, 16, 39, 11, -20, -15, -3, 24, -27, -11, -6, -9, -27, 9, 3, -26, 11, -22, 2, -20, -8, 6, -6, 18, 6, -16, 3, 3, -16, 12, 20, 4, -17, 12, -2, 62, -6, -7, -14, -5, -40, 32, 29, 12, -46, 26, -6, 15, 12, 10, -17, 77, 21, 17, -16, -21, -9, -9, -20, 30, -25, 10, 27, -28, -15, 17, 30, 74, -12, -21, 6, 10, -22, 32, -3, 21, -48, 16, 8, 10, 0, 21, -35, 17, 29, -14, 7, -45, -15, -19, 18, 9, 18, 22, -1, -34, 18, -8, 16, 52, -1, 40, -5, 15, 34, -2, 21, -25, -49, 16, 9, -9, 26, -71, 1),
    (-27, 33, 7, 47, -20, -44, 0, 48, -30, 0, -12, 5, 21, 7, 25, -3, -8, 37, 54, -13, -10, 23, 23, 18, -4, -11, 10, 20, -11, -48, -34, 34, -49, -8, 12, 58, -30, -5, 3, 58, 3, -21, 53, 11, -23, 16, 73, 22, -3, 5, 1, -50, 13, 21, 25, 41, 24, -3, 6, 5, -4, -53, -53, 37, -37, -4, 30, 45, -40, 9, 73, 7, 10, -33, 87, 4, -12, 12, 45, -1, -3, -2, 1, -35, 5, 2, 42, 36, 22, -22, 4, -28, 13, -12, 15, 22, -13, 0, -31, 54, -1, 17, 9, 50, 18, 14, 41, 24, -27, -3, 35, -10, 11, 6, 34, -30, -32, 4, -62, 21, -13, 26, 8, -1, 34, -23, -31, 64, -25, 41, -40, 40, -37, -26, 54, 22, 23, 25, -17, 52, 4, -21, -55, -8, 47, 35, 31, -38, -11, -2, 11, 5, -1, -20, -13, 23, 5, 36, 3, 2, -5, 7, 10, 15, -12, -45, 30, 6, -50, 76, -67, -57, 22, -32, -51, -24, 19, 9, 52, -30, -44, -38, 3, 21, -7, -32, -4, 27, -40, 6, -18, -21, -65, 65, -31, -19, 10, 10, -19, 41, 54, -24, -1, 44, 5, -31, -39, -20, 45, -19, -68, -19, -4, -19, 11, 3, -2, -25, -31, 47, -33, 10, 5, -40, -26, 19, -10, -70, 25, 14, -13, -20, 21, 26, -8, 40, 17, -28, -30, 18, 16, -17, -9, -9, 8, -29, 8, -3, 4, 24, -4, 29, -7, -3, 30, -53, -12, -10, -51, -33, -15, 34, -16, -13, -52, 14, 6, 6, 3, 35, 54, -3, -1, -12, -3, 20, 8, 18, 21, 2, -3, 23, 15, -8, 7, -92, -31, 37, -6),
    (-16, -3, 34, -10, -29, 5, 16, -23, 4, -17, 6, -41, -9, 20, 31, -16, -23, 18, -39, -18, -28, -21, 31, -6, 6, -50, -29, -6, 36, 26, -27, -1, 35, -33, 19, 10, -44, 52, -43, -54, 22, 1, 18, -42, -41, 28, 41, 1, -42, -6, -41, 4, 30, 34, 34, -24, -16, -21, 27, -66, 15, -16, -40, -2, -42, 54, 3, 20, -10, 27, -23, 27, 5, -22, 57, -9, -6, 5, -8, 5, -4, -1, -1, -25, 13, 57, -26, 24, -19, 29, 41, -63, 49, -1, 0, 30, 7, -30, -65, 41, -8, 7, -19, -34, -22, -55, 35, -67, -32, -1, 38, -11, -28, 14, -45, 22, 24, 12, 34, -28, -52, -43, 8, -38, 17, -15, 2, -37, -40, 9, -75, 15, -17, 43, -75, 17, 25, -37, 35, -39, -41, 59, 19, 34, -19, 52, -24, -47, -26, 83, 5, -26, -43, 9, 29, -69, 57, 6, 5, -1, -43, 44, -9, 8, 1, 6, -9, 44, 23, 2, 6, -1, -35, 23, -46, -14, 80, 16, -42, -31, 7, 47, -14, 30, -11, 14, 20, -18, 2, 26, 12, 25, -8, -37, 6, -14, 10, 60, -23, -11, -7, -40, -2, -16, -40, 19, 36, 4, -12, 56, -9, -25, -6, 41, 41, 14, 5, 18, 31, -27, 55, -27, -8, -36, -30, -2, -44, -13, -8, 23, -44, 10, -12, -26, 46, -28, 11, 24, 29, 3, 8, 76, 15, -86, -23, 45, 13, -12, -14, -8, 19, 15, 45, 3, 10, 35, -29, 40, -13, -27, 1, 10, -11, 16, 2, -18, -7, -44, -12, 1, -39, -19, 43, 39, -13, -13, -1, 23, -9, 15, -17, 11, -22, -2, -20, 24, 37, -8, -4),
    (0, -9, -18, -12, -35, -9, -14, -15, -12, -7, 13, -25, -24, 1, -6, 13, 2, 10, 16, -17, 38, 2, 18, -26, 32, -1, 24, -16, 23, -3, 33, -31, -6, -3, -25, -79, -7, 18, 6, -27, -21, -26, -7, -36, -10, 39, 2, 15, -24, 10, 4, -28, 9, -25, -4, -39, 22, 13, 27, -53, 32, -19, 14, -17, -6, 4, 0, -64, 9, -16, -3, 21, 43, -10, -29, -8, -75, -8, 8, 27, -13, 15, -13, 18, 11, -19, 51, -16, -21, 3, -28, -73, 11, 23, 2, -26, 27, -9, 19, 48, -13, 9, -7, 3, -34, -3, 37, 1, 10, 5, -33, 15, -11, -37, -1, -50, 13, 30, -45, 45, -7, 31, 44, 5, 24, -26, -25, 33, 27, -27, -45, 4, -19, 38, -7, -22, -51, -9, 66, -63, 3, 32, 2, 34, -3, -30, -1, -33, 41, 34, -44, -9, 27, 4, 83, -45, 46, -8, 34, -19, -6, -1, -22, -2, 13, -3, -3, -1, 13, -56, 36, -60, -65, 26, -7, 54, 14, 10, 15, -17, 4, -9, -7, -39, 8, -2, -16, -49, 87, 12, 0, -25, 34, -11, 17, -17, -26, -16, -78, -5, -31, 11, -45, -14, 5, 13, -14, -42, 19, -12, 15, 9, 45, 7, -26, 5, 26, -5, -14, -24, 28, 27, 8, -3, 21, 1, 5, 0, -21, 21, -14, -11, -38, 2, 25, -27, 11, 14, 3, -8, -57, 10, -18, 3, 45, 6, -9, 3, 44, 2, 19, -21, 43, 20, 20, -33, 31, 14, -6, 4, 11, 7, 22, -25, -25, -47, 2, -45, 19, -1, 11, 27, -43, 31, -32, -17, 8, -15, 1, -10, 51, 7, 45, -41, 47, -26, -27, -4, -2),
    (17, -1, -17, -24, -18, 42, 8, -12, 16, 44, -25, 10, -3, 6, -23, -9, 29, -1, 20, -34, 6, -30, 9, 12, 41, 34, -6, 10, 29, 17, 9, 14, -4, -33, 17, 10, 10, 3, 30, -54, 7, 12, 1, 33, -31, -15, -41, -6, -19, -9, -7, 10, -2, -21, 1, -13, 53, 9, -25, 46, 2, -24, 9, -20, 36, -17, 42, 22, -20, -6, 15, -61, 13, 32, 0, 34, 15, -2, -37, -11, -34, -6, -3, 66, 25, 17, 0, 8, 33, 11, -16, 27, -21, 11, 7, -13, 30, -3, -34, 13, -20, -30, 39, 14, 23, 13, 30, -24, -28, -4, 44, 14, -31, 19, 67, 23, -30, -22, -5, -11, -13, -28, 6, -17, -19, -47, -1, 24, 5, 28, 13, 24, 25, -40, 34, 30, 4, -12, 61, -25, -52, -8, 67, -16, -31, -29, 45, 27, 7, -43, -31, -39, -23, 6, 1, 21, -72, -60, -34, 29, 3, 13, -4, -5, 12, -39, 35, 2, -14, -37, 9, -55, -18, -26, 46, -16, -1, -25, 37, -8, -37, -20, -59, -48, -5, -8, 11, 38, -47, -42, -34, 14, -10, 14, -3, 0, 36, 10, 24, 21, -20, -14, 59, -7, -1, 36, 59, 8, 28, 16, 13, 4, -21, -14, -38, -19, -3, 17, -6, -3, -6, -31, 1, -19, -61, -7, 2, -3, 35, -19, 42, 52, -9, -46, 40, -16, 18, 57, 48, 21, 57, -5, 3, -74, -27, -4, 10, -15, 18, 27, 15, -23, -1, 2, -28, 42, -61, -5, 26, 1, 19, -15, 21, 37, -39, -32, 56, -18, 1, 35, 12, 0, 60, -2, -6, -79, -2, -7, -31, 2, 16, 49, 24, -4, 1, -31, 5, 25, -12),
    (42, -38, 33, 29, 35, 34, 71, 9, 36, -31, 72, -15, -14, 6, 14, 4, -54, -16, -2, 50, 26, 13, -48, -16, 7, -51, 13, 25, 4, -1, 24, -9, 59, -43, 7, 50, 18, -28, 46, -27, 58, -10, 38, -14, 21, -7, 23, 6, -51, 0, 6, 53, 17, 16, -34, 16, -17, -19, 11, -39, -5, 29, 35, -10, 14, 6, 6, -43, 15, -31, 15, 0, 42, 20, 43, 11, 12, -11, 26, 19, 7, 11, 20, 21, 10, 33, -21, 24, -6, -37, -14, -43, -4, 9, 5, -16, 66, -38, 31, 32, 44, 22, 12, -16, -25, 58, 2, 28, 10, 2, -31, 4, -50, -59, 6, 49, -8, -20, -49, -15, -7, -27, 23, 19, -8, 14, -2, -28, 71, -103, 74, 28, 44, 16, 35, -44, 40, 11, -1, 10, -4, -36, -49, -2, -55, -55, -5, 38, 21, -14, -71, -15, 19, -9, 0, -2, -28, 14, 23, -14, 47, -74, -4, 5, -27, 18, -11, -27, 46, 31, -34, -7, 37, -3, -47, 1, -24, -31, -7, 24, 22, -6, -20, 1, 9, 8, -28, -1, -16, -12, 36, -50, 5, 9, 24, -17, -7, 4, -26, 14, -1, -37, -26, 42, -35, -3, -1, -24, 23, -12, 2, 25, -21, -12, 28, -33, 24, -49, -32, -11, 3, -51, -2, -65, 17, -37, 42, -17, -6, -6, 18, -45, 39, 1, -22, 25, -6, -31, -13, -36, -60, 17, 0, 26, -27, -11, -52, -28, 13, -15, -14, -13, 11, -46, 26, -55, 34, -40, 0, -33, -29, 37, 27, -37, 32, -5, -13, -1, -28, -15, 1, -47, -38, 0, 18, 35, 3, -3, -2, -2, 18, -30, -24, -22, 24, -18, 2, -61, 7),
    (-5, 37, -45, 14, -3, -1, 10, 27, 45, -47, -15, -17, -35, -5, 49, -25, -28, 6, 9, 4, 12, -54, -62, -27, -53, -14, -25, -16, -4, 14, -21, 5, 9, 26, -58, -10, -36, -24, -29, -2, 42, -50, 45, -41, -65, -1, 57, 1, -26, 0, 62, 54, -14, -11, -59, -1, -65, -31, -31, -42, -18, -29, -9, 2, 31, 39, -8, 29, -26, 27, -7, -5, 8, -20, 39, -11, -27, 40, 30, 12, -20, 4, 2, 30, -3, 4, -27, 18, -30, -9, 21, -1, 22, -8, -29, 17, -35, -4, -2, 45, 19, -2, -11, 72, 18, -94, 72, -19, -14, 28, 52, 32, 62, 35, 12, 7, 12, 21, -14, -29, -26, -13, 1, -25, 19, 15, -4, -21, 13, 34, -101, 11, -2, 25, -21, 70, -47, -97, 65, -2, -17, 20, 48, -21, 127, -5, 6, -41, -36, 25, -30, -30, -23, 1, 15, -8, 0, -44, -1, -15, 4, 31, 13, -6, 18, -3, -55, 6, -16, -20, 22, 15, -28, -5, 6, 19, 114, -10, -18, -32, 7, 32, -31, -50, -13, -18, 15, 4, 17, -9, 1, -11, -19, -17, -5, -25, 8, -11, -11, 31, -29, -25, 21, 38, -10, -17, -32, 24, 32, 23, -24, -16, -16, 23, -11, -4, 3, 24, 2, 33, 40, 4, 23, -9, -49, 10, 33, -20, 21, 21, -6, 8, -15, 13, -1, 33, -13, -29, -66, 7, 69, 17, 9, -20, 7, -6, -2, -19, 25, 43, -32, 59, 56, -11, -1, 17, -23, -26, -14, 5, -4, -8, -18, -26, 16, 51, 6, 26, 3, -12, -14, -9, 12, 16, 46, -4, -19, -8, -29, -15, 31, 6, 8, 27, -5, -13, 0, -10, -7),
    (-20, 27, -56, -16, 1, 36, 11, 12, 4, -61, 49, -36, 4, 31, 1, 24, 37, 10, -3, 13, 43, 36, -46, 6, 2, 19, 32, -18, 7, 6, 15, 10, 4, 52, -82, -2, -11, 48, -34, 17, 16, -99, 25, -10, -4, 9, 54, 47, 43, -21, 6, 5, 29, 22, -52, 7, 14, -29, 28, -18, -53, -24, 7, 36, -4, 60, -35, -29, -34, 2, -6, 22, -17, -66, 66, -15, 2, 1, 8, -13, -27, -4, 23, -4, -46, 4, -36, -3, 29, -23, 15, -17, 1, -10, -8, 2, -19, 0, -54, -9, 29, 34, -33, 2, 0, -35, -26, 18, 12, 4, 35, 43, 12, 18, -7, -19, 12, 53, -48, -3, -44, -10, 8, -19, -51, 1, 18, 15, -1, 42, -49, 25, 0, 14, -63, 29, 19, -21, -23, -19, 8, -29, -5, 10, 62, 27, -15, -59, 17, 40, -33, -8, -42, 12, -7, 6, -25, -1, -13, 48, 5, 0, 25, -27, -11, -57, -25, 45, -3, -8, -21, -11, -18, -25, 4, -3, 10, -9, -25, 22, -24, 22, -35, -6, -15, 13, 19, -25, -17, 29, 7, -25, -29, -49, 2, -41, 3, -33, 13, -3, -1, 26, 14, 25, 16, -44, -55, -11, 25, 0, 2, -23, -16, -16, -22, -22, -9, -24, 11, 13, 0, -24, 10, 0, -51, -44, -29, -33, 10, -65, 52, -9, 18, 40, -21, -17, 18, -6, -37, -39, 27, 25, -42, -43, -9, -37, -6, -8, -11, -7, -11, -38, 10, -23, -13, -9, -11, 1, 21, -14, 19, 8, 33, -24, 11, 42, -20, -9, -13, -19, 24, 17, 18, -15, -19, 16, 16, -10, -41, -15, -28, 1, -26, -58, 15, -17, -1, -52, -6),
    (-47, -45, -6, 3, 0, -11, -10, 12, 3, -60, 8, 20, 3, 10, 8, 30, 15, -34, -93, -62, -15, 19, 24, 12, -32, -11, -11, -6, 2, 8, 3, 28, -33, 41, 0, 6, -13, 4, 15, 17, 28, -47, 19, 10, -23, -10, -8, 3, 18, -28, -72, -55, 8, 71, -20, -4, 6, -37, -14, -10, 19, 43, 26, -27, -18, 14, -5, 10, 12, 2, -10, 34, 39, -9, 20, 35, 9, -8, 33, -4, -9, 16, -33, -13, 8, 51, 13, 18, -10, -11, 14, 18, -12, 53, -12, -2, 19, -55, -7, -15, 7, 31, -37, -45, 10, -71, -16, 33, -5, -32, -36, 22, -18, 35, -37, -44, -15, 52, 15, 16, -8, 14, -8, -3, 46, 27, 5, -26, -8, -19, -35, -13, 12, -9, -37, -27, 3, 9, -20, 33, 4, -59, -88, 0, 16, 63, -40, -47, -23, 53, 7, 47, -3, -20, 5, 8, 76, 60, 21, -59, -2, 8, -5, -26, -12, 5, 20, -18, -28, 32, -28, 38, 34, -50, -83, -16, 46, 49, -7, -26, -24, 37, -9, 15, -3, -4, -23, 21, 48, 25, -15, -88, 31, -29, -11, -26, -7, 3, -51, -40, -5, -39, -35, 3, -19, -43, 6, 12, -27, -1, -5, 15, -11, 18, -7, 0, 4, 3, 16, 63, 2, -38, -10, -18, 21, 19, -18, -44, 24, 13, -17, -48, 29, 0, -29, 14, -5, -24, -32, 5, 25, 59, 3, 26, -27, 8, -35, 1, 3, 8, -17, 21, 22, -4, 31, -57, 30, 5, -13, -57, -8, 28, 2, -33, 5, -7, -20, 20, -5, -6, -21, 4, 20, 28, 22, 51, -2, 26, -34, 0, 5, 34, 30, -9, 6, 9, 18, -22, -13),
    (-15, -17, -23, 17, -20, 11, -30, -19, -13, 14, -35, -22, 3, -36, 7, -7, 13, 5, 17, 33, 17, 18, -8, -23, 0, -25, 16, 6, 20, 9, 7, -52, -56, -42, -27, -2, 11, -12, -62, -47, 4, 29, -75, 6, -25, -15, 14, 32, -17, 19, 9, 18, -19, 28, 2, 20, 11, 14, 45, -12, 11, -31, -32, -23, 5, -8, -38, 9, 0, -5, -42, -30, 8, 27, -21, -8, -1, 17, -1, 2, -42, 14, -9, 9, 4, 15, 27, 16, 4, 30, 60, -15, -11, -48, -7, 40, -2, -13, -3, 44, -12, -21, -33, -11, -24, 9, 9, -26, 17, 56, 32, 28, -62, -28, 39, 20, -2, 31, -11, -10, 18, -6, 20, -37, -37, -48, -39, 3, -44, 52, -20, 9, 22, 10, -21, 42, -37, -33, -20, -47, -3, 56, 66, 4, -5, -14, -6, -40, -13, 35, 36, 22, -3, -20, 23, -49, -22, -48, -76, 49, -17, 52, 24, 21, -19, 40, -11, 52, -15, -48, 36, -16, 6, 54, 39, -10, 23, -2, -24, -52, 3, 65, 8, -22, -9, -6, 31, -37, 12, -50, -33, 29, 3, 33, 31, 33, -12, 14, -2, 41, -41, -12, 52, -17, 2, 45, 43, 9, -9, 20, -1, -30, -13, 16, 23, 10, 29, -18, -17, -3, 4, -8, -24, 8, -12, 17, 28, 14, -46, -13, -29, 61, -64, 8, -3, -71, -4, 31, 10, -20, 37, 4, -32, -29, -15, 25, -33, 8, 6, 2, -8, -18, 34, -14, -11, 61, 18, -25, 36, -29, -50, -59, -38, 39, -8, -47, -5, -56, -28, -13, -39, 6, 52, 44, -77, -25, 16, 21, 2, -47, -5, -30, -21, -43, 10, -45, 23, 15, 7),
    (33, 7, 1, 33, -33, 47, -13, -34, 12, -49, -30, 33, -10, 4, -14, 7, -14, 7, -50, 3, -8, 1, -81, 11, 52, 3, 51, 15, -42, 19, -1, -20, 41, -39, -31, 35, 20, 42, -48, 7, 12, -17, -11, 12, -1, 13, -55, 26, -14, 25, -15, -1, 60, 28, -102, -2, 4, 2, 58, 28, 10, 8, 49, -52, 12, -43, -51, 21, -8, 4, -44, -29, 18, -18, 8, 11, -28, -24, -33, 2, -12, 42, 8, 12, -2, 4, -87, 5, -15, 38, 56, 4, -3, 7, 55, -32, 28, 9, 35, -63, -13, 47, -72, -15, -66, -8, -51, -5, 10, -12, -22, -18, -4, 82, -5, -21, -9, 1, -45, -6, 11, -45, 31, 15, 2, -8, -23, -56, 70, -57, -19, -42, -17, 24, -57, -75, -48, 22, -39, -37, 7, -5, 12, -17, -14, 46, 0, -2, 9, 21, 7, -29, 17, 8, 26, -29, -44, 22, -20, -84, 48, -68, 20, 4, 14, 35, -53, -36, -45, -3, -22, -31, -4, -20, -4, -17, 24, 27, -11, 10, -22, 13, 30, -21, 30, 23, 47, -50, -32, -48, -9, -22, -15, -27, 54, -25, -21, -7, -10, -33, 12, -43, 8, 14, 7, -10, 4, -35, -4, 54, 9, 9, -36, -14, 26, 4, 7, 6, 25, -28, 22, 22, 21, -28, 29, -21, 49, -48, -11, -12, -7, -11, 4, 18, 21, 17, -26, -19, -2, -2, 21, 41, -15, -31, -16, -26, -25, 15, 5, 6, -12, 10, 29, 31, -1, -56, 4, 28, 43, -43, 30, -11, 14, 23, 8, 32, 12, 16, -10, 19, 6, -8, 34, -21, 5, -47, -42, -6, 15, -15, -10, 41, -44, 23, 46, 37, 29, 8, -5),
    (-14, 44, 8, -16, -31, -14, -7, 34, 6, -50, 40, 4, 7, 11, 32, 52, 45, -27, -14, -2, -39, -5, -35, -5, -44, -38, -29, -16, -19, -16, -12, -8, -37, 93, -30, -40, -9, 0, -23, 46, 38, -36, 58, 19, -24, 32, 64, 14, -21, 5, -3, 18, -31, 18, 0, -6, -59, -15, -9, -29, 15, 2, -23, -52, 1, -2, 8, -19, -13, -16, -26, -6, 31, 12, 33, -7, -20, -7, 62, 5, -51, 42, 19, 51, -9, -12, 26, 4, -13, -45, -17, 0, 11, -12, -36, -92, 11, 53, -74, 30, -16, 38, -4, 54, 16, -7, 41, -8, -24, 1, 67, -16, 51, 31, 14, 13, 23, 20, -10, -4, -54, -35, -7, 29, -25, 25, -10, 15, 26, 16, -42, 2, -22, 16, -60, 43, 33, -31, 60, -23, -42, 0, 94, -20, 44, 4, -25, 35, 25, 58, -34, -49, -82, -44, 1, -10, -46, 2, -27, -21, -12, 36, -17, 13, -26, 47, -55, -10, 38, -35, 41, 1, -31, 24, 42, 15, -12, 25, 39, 41, -30, 42, -32, -33, -72, 5, 9, -27, 10, -17, -48, 2, 16, 3, -33, -40, -4, 6, 21, 48, 9, -15, -15, 24, -3, -14, 23, 26, 27, 10, 27, 18, 7, 22, 6, -28, -48, -9, -10, 23, -29, 15, -9, 4, 27, 26, -41, -15, 3, 48, -24, 37, 10, -49, 14, 0, -48, -6, 53, -1, 39, 38, 34, 30, 27, 60, -16, -15, -88, -3, -14, 5, -26, 16, -6, -35, 1, 50, -28, -13, -6, 31, -3, 37, -1, -4, 17, -8, -17, 31, -9, -17, 42, 33, 14, 23, 0, 43, 17, -19, -34, 7, -21, 26, -24, 13, -6, 7, 8),
    (0, -21, 31, 23, -21, 1, 1, -31, 15, 26, 7, 17, -21, -35, -14, -10, 0, -19, -36, -1, -16, -16, 19, 16, -14, -4, -21, 18, 9, -5, -24, -10, -1, -32, 40, -16, 14, 5, -13, 1, 10, 33, 26, 49, 16, -41, 27, -1, 3, 7, -29, 9, -15, -9, -10, 36, -35, 10, -33, 22, -9, 56, 14, -34, -12, 12, 6, -14, 12, 3, 17, -6, 16, 63, 12, 19, 7, -57, 11, -41, 14, 15, -7, -17, 10, 5, 22, 63, -36, -34, -20, 47, -3, 45, 4, -34, -6, -12, 14, 36, 21, 1, -9, -66, 34, 10, -52, 40, -20, -19, -56, -14, -18, 23, 2, 26, -12, -8, -26, -8, -60, 10, -29, 35, -52, -12, -50, -26, -1, 29, -43, -47, -14, -33, 24, -68, 38, 11, -74, 98, 20, -61, -47, 3, 13, 22, 20, 41, 3, -14, -23, -9, -68, 19, -11, 85, -67, 15, -8, -84, -35, -15, -4, -9, -7, 18, 12, -42, 14, 29, -43, 51, 37, -27, -22, -10, -13, -43, 14, -1, 7, -4, 12, 18, -8, 8, 22, 46, -23, 8, -4, -55, -4, 17, -7, -31, 21, -5, 24, -52, 19, 3, -10, 66, -5, -10, 0, -1, 7, 28, 13, 32, -22, 31, -52, -21, -8, 1, -17, 53, -19, -31, -18, 22, 34, 42, -32, 25, -40, -16, 43, -18, 25, 4, -48, 48, 27, -6, -21, 18, 30, 39, 46, -10, 3, 6, -44, 23, -7, -15, -25, 38, -51, 24, 3, -5, -8, -12, -14, 1, -13, 2, 9, -2, -1, 17, -24, 2, 35, 32, 13, 34, 5, 12, -4, -9, 3, 9, 5, 1, -3, -2, -15, 22, -21, 6, -10, -16, -4),
    (0, -52, -4, 8, -58, 4, -17, -34, 23, -20, 4, 20, -3, -48, -39, -9, -44, -16, -4, -7, 30, 14, 49, -3, 19, -5, -16, 27, 12, -19, 44, -24, 71, -13, 19, 30, -47, 41, 23, -17, 26, 27, -8, -13, 3, -44, 21, -13, -80, -8, 62, 68, 54, 49, 1, -5, -33, 0, 2, 4, -18, 5, -2, -9, 55, 26, 5, -42, 16, 35, 3, 29, 18, 11, 22, -23, -26, 2, 40, -44, -12, -12, 53, 73, 14, 7, 6, -26, -20, -54, -27, -8, -48, 7, 16, -6, 51, -47, 8, 20, -39, -16, -35, 4, 6, 2, -50, 13, -17, -10, -8, -1, 1, 7, -28, 12, -10, -3, 69, 4, -30, -18, 10, 0, 19, 44, 25, -21, 57, 11, 34, 7, -23, 29, -13, 23, 26, 15, -12, -33, -20, -19, 80, -16, -28, -35, 23, 24, -3, 29, 3, -30, -66, -55, -7, -67, -7, 47, 5, -18, -5, 63, 30, -5, -18, 28, 4, 47, 13, -10, 27, -36, -12, 12, 32, -13, -8, 10, 0, 39, 44, 47, -3, -6, -80, -39, -2, -45, -24, 38, -20, 10, 30, -20, 58, -9, -7, 36, 2, 23, 5, 32, 7, -9, 29, -16, 2, -35, 0, -10, -24, 46, -16, 6, 18, -18, -35, -10, -3, -6, 24, -6, -2, -58, 21, 16, 17, -3, -12, 4, -89, 41, -6, -18, 27, -50, -12, 15, 54, 6, 4, 27, -10, 32, 18, 1, -6, -27, -32, -12, -16, -57, 21, -8, 21, -19, -33, 40, -21, 11, 8, 24, 26, 37, 12, -1, 0, -31, 19, 7, 27, 10, 82, -5, -28, 0, 2, 23, 6, 11, 12, -1, -1, -41, 11, 16, 33, 18, 11),
    (-12, 5, 40, 19, 27, -1, 0, -33, -29, 1, -64, -25, 28, 32, -60, -9, 28, 0, -28, -25, -4, 10, 40, 14, 9, 2, -21, -10, 69, 33, 14, 11, -55, 20, 14, 18, -3, -8, -19, -31, -40, -21, -24, -6, -8, 37, -91, 57, 41, -2, -55, -2, -2, 14, 77, 19, 19, 29, -2, 2, 97, 19, 17, 21, -36, 5, 5, -8, -13, -21, 10, -19, -30, -44, 10, 3, 3, 6, -71, 10, -6, -1, -39, -4, -13, 20, 5, 7, 34, -38, 3, 34, 14, 11, 13, 7, -5, 1, -11, -22, -4, 20, -13, -31, -46, 27, -16, -7, 37, 26, -31, 4, 12, 0, -10, -3, 45, 38, -1, 17, 12, 9, 28, -32, 15, 4, 15, 9, -6, -23, -66, 21, 24, 43, -13, -53, -26, -50, -24, 9, -14, 32, -74, 28, -26, 13, -1, -37, 45, 29, -27, 28, 62, 14, 15, -11, 76, -26, -1, 48, 34, -37, -34, 25, -35, 6, 6, -66, -38, -24, -20, -10, 26, 10, -62, 21, -60, 1, -8, 8, 22, -2, 37, -18, 68, 16, 16, -4, 13, -29, 9, 26, 20, -15, -5, -5, 3, 3, -45, -24, -41, 20, 21, -35, 21, -1, 9, -16, -11, -8, 1, -33, 6, -3, 27, -12, 21, -3, 21, -36, -21, -46, 13, 7, -14, -39, 18, -2, 3, 6, 8, -21, 14, -40, -24, -12, -16, 21, 4, 32, -66, 29, -9, -41, -6, 41, -11, 44, 48, 10, 23, 6, -39, -10, -13, 5, 32, 1, -1, -2, 19, 21, -19, 2, -18, -26, 12, -43, -43, 28, 11, -6, -33, 2, -18, -4, -9, 6, -41, 25, 8, -38, 13, 23, -11, -14, -46, 21, -6),
    (5, -11, 13, -37, 19, 20, -31, -19, -5, 8, -12, 7, 3, -47, -17, -21, 29, -44, 2, -54, 8, 16, -60, 6, 38, 24, 37, 54, -44, -14, 29, -36, -4, 13, -17, -15, 6, -15, -52, -28, -20, -23, -8, 10, 27, -19, 19, 21, 31, 18, 0, -67, -30, 48, -65, -20, -5, 3, 10, 41, -32, -49, 14, -28, -20, 30, -38, 0, 15, 18, -38, -14, -33, 18, -19, -15, 23, 2, 26, -12, 33, 39, 10, -23, 6, 32, -9, -16, -24, 20, 3, 2, -17, -31, 14, -13, -39, 50, -2, -61, -2, 25, 43, 4, 23, -40, -13, 47, 33, -43, 9, -1, 55, 50, 10, -55, 38, 6, -32, -27, 7, -8, -22, 65, -70, -5, 9, -40, -52, 58, 12, -67, -11, 8, -14, -13, -41, -32, -15, 77, 42, -52, 34, 0, 67, 53, 12, -76, 12, -16, -25, 5, -14, 36, -15, 93, -75, -15, 8, -56, -42, -1, -10, -30, -8, -19, -36, -2, -47, -22, 11, 16, 26, -17, 19, 24, 59, 24, -5, -39, -22, -6, 27, 10, -20, 13, -14, 48, -43, -12, 10, -20, 16, 20, 36, -1, -13, 8, 28, -2, 5, -2, 9, -9, 10, -12, -37, 18, 44, -31, 32, -40, 2, -8, -50, -26, -27, 13, 16, 16, 9, 10, 15, 11, 27, 25, 4, -18, -33, 7, 10, -7, 8, -63, -31, 77, 16, -27, -37, 34, 3, 14, -19, -23, 14, -20, -7, 12, -31, -8, -15, 57, -32, -5, 9, -17, 6, -18, -24, 2, -11, 11, 1, 14, -7, -62, 1, 24, -6, -13, -35, 42, 11, 32, -3, -21, 4, -4, 6, 32, -28, 22, -11, 21, -7, -28, 1, -27, -8),
    (-20, 1, 41, -28, -40, 14, 5, -61, 37, 10, -16, 40, -35, -38, 46, -7, -14, -53, -8, -33, -5, -18, 11, 17, -16, -32, 10, -12, -26, 12, 21, -26, 22, 14, 6, 2, -13, 12, -9, -13, 36, 50, 24, 31, -22, -24, 38, -37, 3, -39, 67, 44, 45, 22, -52, -8, -41, -36, -30, 41, -48, 30, -12, -29, -7, 13, -22, 11, -16, -24, 10, 30, 24, 2, 7, -5, -9, 1, 1, 2, -2, -18, 30, 37, -20, 33, -4, 17, -27, 13, -12, 16, -21, 16, -28, -13, 31, -22, 52, 20, -37, 21, 29, -14, 14, 95, 7, 3, -49, -39, 10, -21, -28, -21, 20, 51, 9, 19, -22, 19, -88, -24, -42, 2, -41, -3, -30, -13, -2, 20, 11, 35, -44, -20, 11, 30, 17, 58, -4, -21, 14, -18, 46, -29, -36, -23, 69, 49, 20, 40, -40, 28, -73, -41, 13, -11, -42, -5, -33, -6, -14, -17, 22, -5, -18, 3, -8, 22, -12, 15, -19, -61, 10, 14, 20, -2, 7, 4, 29, 26, 33, 49, -28, 33, -21, -7, -3, -31, -13, -10, -42, 4, 25, -27, 9, 42, -15, 40, -33, -11, -9, 24, -17, -15, -7, -20, 54, -29, -36, -6, 15, 50, -17, -10, -36, 10, -67, -13, -16, 16, -26, 5, -32, -16, 1, 19, 32, 41, -13, 4, 26, 28, -7, 52, 7, -67, 13, 34, 79, 6, 12, 17, 38, 31, 28, 27, -25, 14, -29, -31, 13, -38, -10, 0, -17, 57, 8, 12, 7, 37, -9, 37, 26, 21, -50, 20, 6, -34, -2, 38, 30, -24, 22, -13, 24, 0, 30, 4, -18, -3, 29, -26, 5, -26, -6, 0, -21, 50, 13),
    (-16, -48, -5, 41, -5, -35, 26, -28, -2, 21, -4, -11, 1, -26, -17, 1, -36, 6, 25, -2, -5, -7, 27, 29, 34, 31, 21, 59, -18, -6, -21, 47, 61, -54, 30, 49, 24, -29, -24, -25, -41, -38, -21, -12, -8, 10, 42, 22, -80, -12, 15, 7, -8, 16, 23, 3, -11, -11, 30, 14, -39, -61, -38, 41, 20, 7, -8, 12, -9, 18, -10, 12, 72, -34, 58, 36, 5, 40, 13, -34, -19, 1, 22, 9, -32, 20, 24, 9, -51, 18, -1, 30, -7, -13, 9, -19, -2, -30, 6, 30, 17, -23, -9, -15, -52, -23, 21, -12, -24, 46, 10, -21, -58, 15, -28, -30, -10, 3, 30, 45, 35, 31, 37, -2, -33, -61, -46, 35, 20, -31, 3, 61, 23, -14, -19, 9, 35, -66, 54, -9, -42, 29, 41, -1, -58, -19, -28, -17, 6, 8, -26, 23, -53, -13, 3, -11, 0, -28, -95, 37, -41, -19, 23, -41, 8, -34, 32, 35, 26, -9, -12, 12, 4, -18, 1, 14, -11, 7, -33, -54, -6, 27, -4, 3, -15, -10, 3, 22, 0, 52, -28, 33, 26, -6, -3, -4, 9, 6, -41, -15, -32, -27, 1, 37, -5, 10, -20, -27, -11, 18, -21, 15, 2, 37, -16, 18, -22, 44, 10, -37, -37, -39, -33, 25, 8, 19, -26, -12, -25, -12, -12, 13, 66, -15, 18, 31, -27, -58, -20, -11, -18, 41, 21, -22, 20, 9, 8, 16, -86, 10, 11, 58, -9, 2, -25, -36, -32, -13, -40, -27, -26, -11, 18, -7, -3, 43, -44, -22, 30, -13, -18, 28, 14, 4, 16, -26, -20, -8, 21, 16, -2, -6, -3, 19, 14, 34, 1, 2, -4),
    (-7, 25, 21, -6, -2, 10, 55, 32, -5, -2, 54, -20, -32, 4, 18, 2, 90, -49, -27, -58, 11, -29, -2, -22, 34, 19, -4, -59, 15, -2, 8, 60, -2, 23, 28, 18, -47, 28, 47, 23, -1, -55, 31, -7, -45, 36, 11, 3, 36, -34, 9, 2, -16, 8, -9, -37, 68, 33, 8, -28, 7, 25, 0, 13, -1, 29, 44, 25, -14, 0, -6, -5, -6, -41, 12, -8, -36, 21, -28, 4, -11, 5, -7, 14, -15, -13, -7, 4, 28, -10, -21, 17, 28, 16, 18, -23, -1, 18, -55, -5, -27, -13, 27, -14, 69, 44, 27, 37, 23, -26, -17, 36, 15, -23, -33, -30, 19, -22, 53, 18, -26, -9, 5, -3, 24, 7, 17, -22, 31, -25, -38, 11, 5, -12, 55, -8, 77, 8, 40, 49, 24, -59, -3, -17, 27, -5, -42, -26, 33, -7, 25, 28, -6, -33, 2, 3, 30, -13, 7, -1, 9, -16, -40, -66, 30, 16, 31, 9, 23, 20, 4, -8, 16, -17, 18, -4, 23, -22, -3, -22, -11, -21, 15, 34, -28, 19, -2, -30, 11, -14, 16, -63, 1, 11, 19, 29, 6, -14, -23, -31, 5, 34, -8, 23, -10, -6, 9, -14, 2, -8, -7, -16, -34, -10, -9, 13, -31, 3, -16, -7, 16, 13, -9, -11, -2, -25, 8, 37, 25, -21, -14, 7, 7, 36, -31, 30, 4, 15, -54, -8, -16, 25, 17, -8, -58, -14, 2, 53, -43, -34, -27, -12, -11, -17, -41, -48, 5, 3, -24, 75, 27, -65, -46, -7, 36, 49, -1, -2, 26, -21, -34, 10, -38, -33, -3, 20, -42, -17, -16, 21, -3, 18, -6, 21, -23, -9, -43, -27, -3),
    (-17, 2, 16, -25, 5, 31, -23, 28, -26, 5, -17, -19, -42, 22, 10, -9, 8, -66, 7, -36, -31, 6, 9, -54, 27, 0, -9, 3, 12, -31, 23, 29, -30, 41, 39, -39, 15, 34, -15, -2, -33, -8, 15, -7, -17, 17, 50, -12, 29, 31, 3, 0, 1, 19, -3, -60, 10, 30, -8, 42, 35, 50, 18, -12, 4, 27, 7, -47, 10, 20, -18, -7, -33, 2, -24, -19, -2, -30, 25, -1, 25, 19, 19, 1, -9, -3, 18, -38, 17, 15, -10, 37, -8, 28, -7, -55, 3, 20, 48, 6, -26, -11, 17, 28, -46, 40, 17, -33, 16, 26, 28, 3, 20, -36, -14, -35, -18, -57, 34, -60, 31, 0, -8, 9, -6, 15, 27, 64, -19, 51, 65, -50, -16, 9, 20, 46, -25, -2, -2, -25, -20, 21, 22, -23, 73, -39, -43, 35, -8, 1, -20, -106, 66, -3, -3, 3, 59, -8, 42, -18, -33, 47, 54, -89, -12, 28, 21, 44, -41, -14, -7, 1, -52, 16, 5, -14, 47, 35, -21, 41, -2, -1, 18, -58, 48, 8, -9, 19, 50, 0, 38, -34, 39, -16, 0, 20, 8, 13, 11, -15, 8, 46, -21, 21, 8, -28, 27, 41, -23, -16, -7, -17, -35, 15, -22, 11, 20, -20, -8, -1, -10, 36, -38, -5, -11, 9, 28, 16, 18, -8, 27, 17, -5, 47, 27, -4, 23, -2, 7, -38, 27, -63, -39, -26, -11, -14, 35, -22, 9, -46, -23, -38, 21, 30, 1, 10, 18, 20, 19, 6, 27, 2, -3, 44, -28, 30, 4, -22, 8, 1, 18, -43, 53, -47, -48, 26, 17, -21, 30, -56, 23, -25, 13, -20, 5, 6, 3, 15, 21),
    (-41, -12, -20, 22, -26, -2, 24, -10, 43, 44, 13, 33, 38, -41, -68, 19, 9, 19, -36, -3, -16, -9, 24, 58, 11, -36, -42, -15, 39, 50, 30, 20, -29, -53, -3, 49, 15, -29, 31, -46, 23, 63, 24, 29, 64, -33, -77, 10, -16, -2, -9, 15, -39, 0, -6, 61, 4, -5, -20, 8, 27, 25, 8, 28, -26, -34, 14, 22, 9, 2, -16, -40, 6, 21, -30, 17, 32, -5, -53, 9, -31, 16, 7, 33, -16, -9, 37, 15, 12, 15, -20, 12, 44, -5, 6, -13, -16, -38, 40, 16, 9, -28, 19, -49, 40, 25, -32, 31, 28, -7, -56, -24, -66, 47, 36, 7, -3, -8, -31, 30, 0, 0, -8, 9, 5, 24, 36, -14, 26, -75, 27, 26, 32, -31, 3, -71, 18, 46, -35, 50, 41, -29, -86, 3, -115, -12, 57, 28, -14, -29, -39, 37, 0, -8, -38, 27, -19, 6, 10, -27, 40, -48, -5, -21, 16, 16, -24, -42, -3, 21, -34, 15, 16, -20, -40, 18, -74, -26, 38, 48, 4, -17, -46, -14, 23, 14, -21, 26, 22, -8, -11, -23, -33, 8, 70, -13, 33, -6, 24, -15, 27, 6, -28, 11, 4, -10, -44, 3, -29, 8, 38, -1, -13, -8, -46, -3, 9, 32, -11, 4, 25, 29, 2, -7, -13, -6, 40, -24, 23, 18, -15, -34, 23, -10, -56, 13, -41, -19, -28, -4, -52, -17, 53, 31, -29, -17, -39, 1, 18, -3, -10, 20, 2, -9, -12, -51, 19, 10, 12, -40, -19, 7, -17, -7, 21, 14, -20, 7, 15, 4, -20, 18, 1, -2, 38, 20, -2, -13, -24, -24, -25, -1, 9, -2, -29, -40, 9, -40, -8),
    (-36, -65, 52, 35, -2, -31, 69, -11, -9, 48, -10, -13, 36, -42, -12, 10, 10, 41, -1, 21, -22, -21, 6, 22, 9, -20, -47, 35, -6, 34, 6, 7, -14, -56, 69, -1, -12, -21, 31, -3, -12, -4, -50, -26, -16, -28, 37, 3, -12, -46, 21, 43, -14, -28, 6, 29, -15, -23, -13, -17, 11, 15, -6, -69, -3, -41, 19, 24, 31, -3, -3, -28, -11, -3, -28, -10, -1, -3, 47, -43, -44, -50, 54, 12, 18, -3, -13, 5, -23, 0, 12, -34, -33, -17, 5, 11, 16, -43, 33, 33, -12, -27, 9, -69, 9, 39, -5, 35, 6, -21, -4, 16, -48, 11, 68, 75, -18, 10, 16, 58, 20, -15, -29, 33, -9, 62, 17, -14, 14, -49, 58, 27, -17, -11, 27, -28, -35, 86, -52, -42, 29, -18, 33, -23, -11, -17, 52, 22, -16, -10, 71, 4, -3, -30, -16, -7, 22, -22, -19, 8, 20, 2, -8, 8, 27, -10, 17, 1, -43, -15, -45, -48, 25, 9, 45, -49, 19, 4, 27, 12, 22, -23, -40, -28, 7, 13, -12, -53, -24, -9, 25, 18, 28, -25, 26, -21, -9, -9, 27, -12, 21, 34, -32, 36, 18, -2, -12, -10, -16, 4, 66, 27, 3, -1, -30, 33, 35, 15, -13, 68, -31, -16, 7, -48, 23, -12, 19, -13, -4, 41, -11, -36, -19, 49, -43, -2, 3, -7, 26, -11, -57, -18, 48, 20, 11, 13, 11, -24, 33, 17, -21, 6, -27, -40, -24, 42, 2, 17, 13, 24, -16, 25, -30, 7, 7, -43, 48, 31, -38, -3, -26, -43, 14, 24, -17, -5, -4, 11, -26, -1, 41, -25, -21, 9, 16, -1, 27, 10, 6),
    (-17, -30, -32, 16, -16, -29, -18, 20, 5, -50, -9, 11, -54, -2, 89, -38, 56, -7, -32, -29, 8, -39, 63, 5, -6, -43, -6, -1, 30, -54, 4, -26, -39, -27, 7, -14, -7, -38, 11, 50, 33, -76, 10, -1, -20, -16, 71, -9, 84, -45, -24, -9, -28, -15, 31, -14, -55, -32, 33, -13, -2, -18, 2, -19, -25, -26, 50, -44, -43, -10, 30, 25, 34, -1, 18, -3, -34, -30, 26, -23, 50, -63, -30, -1, 8, -8, 35, -25, -38, -15, -23, -54, -19, -5, -38, -41, 11, -56, -6, 34, -26, 40, 47, 29, -10, -7, 29, -49, 17, 38, 48, -8, -1, -22, -5, 9, 36, 12, 0, -21, 21, 1, 31, -28, 36, 3, -18, 10, -7, 31, -44, 39, 24, -17, 52, 42, 19, -46, 26, -37, -9, 43, 81, 19, 48, 55, 3, -16, 21, 9, -20, -26, 3, -33, -5, -38, 39, 11, -21, 29, -20, 11, -5, 33, -15, -5, 34, 25, 13, -8, 14, -13, -29, 45, 70, 29, 23, 46, 17, -21, -22, 22, -8, 7, -37, 7, 13, -39, 11, -1, -21, -42, 28, -37, 52, 20, 9, 25, 2, 15, -37, 17, 27, -70, -4, 21, 47, -13, -7, 25, 23, 16, 7, -12, -6, 13, 0, -20, 10, -22, -10, 13, 1, 13, 13, 5, 4, 11, -19, 10, 5, -9, 16, 1, 59, -27, -5, -5, 71, 11, 26, -12, -6, 36, 11, 11, 3, 0, 17, 12, -17, -32, 28, 20, 22, 33, 27, 22, 0, 1, -38, 9, -9, -6, -3, -12, 49, 14, -14, 8, 60, 4, 22, -28, -14, 27, 36, 12, 0, 10, 4, 9, -5, -1, -3, 15, -6, -14, 14),
    (-48, 7, -34, 1, -33, 9, 22, 38, 29, -12, 22, 67, -23, 20, -7, 0, 28, -1, -42, 3, -17, -30, -35, 0, 16, -23, 29, -25, 45, -12, -30, 23, -29, -21, -22, 24, -55, 22, 39, -40, 13, 28, -39, 76, 27, -34, -77, -20, 12, 4, -29, -8, 22, -9, 22, 32, 7, 13, 24, 36, -22, 25, 51, -3, 26, -30, -15, 26, 26, 13, -13, -48, -39, 22, -45, 32, -7, -13, -40, -26, -24, -2, -13, 38, -29, 4, -2, 32, 11, -7, -4, 44, 1, 0, 28, 28, -33, 43, -18, -34, -4, 35, 8, -4, 47, 13, -35, 84, -24, -36, -63, 10, 54, 33, -15, 37, 34, -18, 1, 15, 31, 5, 6, 40, -10, -1, 24, -12, 79, -60, -50, 35, -21, -4, -3, -65, 25, 58, -93, 97, 28, -8, -75, 11, -59, -45, -7, 12, 47, -23, 14, 20, 21, 2, 11, 81, -60, -34, -11, -18, 61, -19, -34, -21, -23, -8, -22, -8, 11, 21, -54, -2, 10, 34, 35, -2, -49, -42, 1, 33, -51, 32, 80, 4, -12, -19, 13, 13, -6, -52, -9, 32, 0, 36, -11, -37, -43, 10, -16, -22, 46, 35, -10, 15, 11, -39, -34, 9, 13, -11, -36, -19, 12, -24, 38, 7, 9, 8, 2, 21, 5, -10, 27, -41, 48, -58, -34, 11, 16, -33, 28, -25, 34, 54, -66, 1, 40, 16, 7, -11, -46, -5, -13, -45, -24, 0, 21, 32, -20, -2, -22, -11, -10, -1, -3, 32, 5, -7, -23, 34, -7, -5, -7, 32, -29, 20, -6, -59, -21, 41, -5, -1, -27, -20, -13, -13, -10, 45, -14, -2, -41, -15, -26, -30, 19, -19, -37, 35, -5),
    (-19, 5, -30, 3, -16, -8, -8, 53, -9, -34, 11, -64, -5, -1, 18, 28, 23, 34, -20, -43, -13, 26, 32, -22, -20, -19, 4, -32, 14, 44, -2, 32, -39, 17, 38, 25, -27, 0, -33, 36, 10, -39, 0, -36, -7, 5, 27, -6, 38, -13, -7, 2, -31, -19, 35, -9, 22, -15, 4, -22, 45, -16, 11, -1, 5, 38, 33, 5, 4, 7, 20, -7, 27, -69, 35, -9, -43, 46, -3, 62, 30, -49, -53, 25, 6, 10, 8, 5, 14, 10, 24, -37, 25, -9, -21, -38, 7, -42, -7, -19, -30, -19, -46, -2, -28, 6, -27, -12, 11, -13, 41, 14, 48, 48, -35, 21, -7, -6, 18, -48, -7, 10, -2, -42, -7, 21, -16, -27, -16, -3, -25, 7, -27, -17, -43, 40, -12, -12, 3, -38, -19, 39, 27, -9, 28, -39, -58, 18, -2, 23, 58, 15, -24, -35, 47, -104, 56, -32, -42, -6, -54, 34, -16, -23, 21, -4, 15, 28, 4, 21, -10, -5, -13, 11, -25, 52, 47, 2, -36, -53, 17, 20, 3, -1, 56, -18, 41, -35, 89, 30, -9, 6, 41, 12, -87, 11, 19, -12, 2, -4, -26, -32, 22, -7, 3, 15, 36, 43, -2, 24, 9, 2, -24, -25, -14, -16, 9, -35, 57, -46, 26, -48, 20, -11, -2, 18, -12, 1, -24, -6, 0, 25, -29, -34, 33, -5, -25, 54, 36, 24, 20, -18, -13, -27, -1, 22, 12, 39, 14, 28, 27, -56, 43, 13, 19, 5, -32, 34, -19, 18, 0, 33, 26, 8, 11, 48, 29, -13, 13, 1, -5, 33, 30, 33, 18, 13, -25, 0, -15, 8, 19, -17, -29, 7, 21, 1, 22, 14, -4),
    (13, 14, -40, 2, -4, -3, 15, -40, 49, 10, -14, 24, 60, -37, -66, -37, 4, 47, -42, -5, 46, -2, -7, 34, 33, -15, -1, -35, -18, 38, 23, -41, -29, -45, -6, 1, 4, 18, 53, -3, 13, 25, 6, 5, 26, -25, -59, 11, 26, 12, -19, -33, 37, 33, 53, 20, 3, 23, 13, -19, 19, 32, 23, -14, -30, -66, 3, -13, -14, -19, 3, 9, -8, 14, -1, 5, -9, 5, 16, -12, 16, 4, -8, -17, 47, -15, 62, -2, -9, 2, 1, 13, -7, 0, 18, -24, 31, -14, 38, -37, -8, -13, -10, -19, 19, 10, -3, -35, 1, -3, 9, 18, 3, 61, 15, 32, 17, 19, -28, -6, -14, -3, 25, -20, 18, 54, -7, -56, 24, -53, 38, -7, 34, -30, -22, -21, 67, 73, -55, -21, -12, -21, 16, 32, -42, 42, -14, 33, 14, -6, -17, 28, -35, -20, -15, -62, 38, 73, 34, -76, -43, -43, 6, 43, 39, -28, -24, 16, 4, 57, -40, -4, 3, -26, 27, -24, -34, 16, -25, -24, -21, 33, 14, 23, 0, -26, 10, -12, 17, 32, -16, -53, 21, -25, 12, 0, -8, -6, -9, 11, -4, -1, 17, 33, -11, 0, -26, -13, -31, -25, 15, 17, -53, -43, 2, -42, -8, 21, -3, 2, 10, -49, -16, -18, 20, -32, 51, -30, 19, 10, -10, -4, 4, 16, -14, 49, -36, -1, -20, -44, -44, 31, 23, 30, -27, -42, -15, -15, 10, 35, -29, 0, 28, -22, 33, -44, 16, 2, 28, 2, 27, 26, 2, -20, -9, -9, -35, 4, -52, 4, 11, -37, -54, 45, 10, 29, -50, 3, 19, 1, 20, -14, -21, 3, 20, -78, -3, 12, 6)
  );
  ----------------
  CONSTANT Flatten_1_Columns : NATURAL := 4;
  CONSTANT Flatten_1_Rows    : NATURAL := 4;
  CONSTANT Flatten_1_Values  : NATURAL := 48;
  ----------------
  CONSTANT NN_Layer_1_Activation : Activation_T := relu;
  CONSTANT NN_Layer_1_Inputs     : NATURAL := 768;
  CONSTANT NN_Layer_1_Outputs    : NATURAL := 10;
  CONSTANT NN_Layer_1_Out_Offset : INTEGER := 4;
  CONSTANT NN_Layer_1_Offset     : INTEGER := 0;
  CONSTANT NN_Layer_1 : CNN_Weights_T(0 to NN_Layer_1_Outputs-1, 0 to NN_Layer_1_Inputs) :=
  (
    (2, -20, -22, 7, 15, -8, -3, 2, 11, -1, -22, -9, -2, -8, 5, -31, -8, -40, -38, -13, -17, -17, 7, -41, 4, 5, -24, -3, 0, 9, -22, 29, 3, -3, -15, 16, -1, -18, -3, 5, 14, 2, -6, -12, 11, -40, 15, 24, 8, -24, -18, 18, 13, 31, -4, 8, -5, 4, -4, -42, 28, -7, 21, -32, 13, -32, -25, 2, -34, -13, 2, -18, -1, 0, -3, 28, -8, 0, -12, -2, 0, -12, -6, 15, -2, -11, 4, -2, 23, 14, 28, 8, 2, -20, 17, 35, 5, -35, -5, 11, 33, 22, -16, 12, -12, -6, 5, -28, 8, -7, 14, -18, 5, 12, -24, 5, -20, -9, -4, -12, -18, 17, 2, 35, -1, 0, 2, -21, -8, -23, -1, -7, 12, -26, 10, -5, 15, 21, 23, 9, 9, -5, 8, 15, 1, 14, 8, -10, 5, 1, -5, -4, 6, 3, 14, -15, 4, -4, 18, -26, -10, -4, 3, -3, -17, 0, -1, -10, 6, -12, -1, -2, -4, -18, 3, 0, -2, -14, 10, 2, 18, -23, 5, -16, 10, 15, 10, 9, 12, -1, 4, 1, -4, -19, -29, 8, 11, 30, -17, -11, 9, 28, 16, -29, 20, -16, 3, -45, -24, -35, -47, 8, 14, 0, 23, -25, 21, -19, -16, 1, 4, 11, -2, 21, 4, 20, -30, -1, -17, -27, 12, 3, 10, 26, 0, 7, 16, -41, 11, 29, 8, -19, -34, 2, 15, 52, -18, -3, 9, 11, 27, -36, 26, -16, 51, -43, -50, -45, -24, -5, -25, 12, 8, -22, 34, -17, -11, 3, -15, -18, 5, 4, -7, -20, -10, -9, -29, -20, 4, -3, 31, 56, 22, 34, 17, -51, 28, 27, 5, -25, -38, 5, 11, 30, 3, 3, -11, -7, 15, 8, 16, -2, 35, -23, -32, -34, -21, 8, -30, 17, 7, -38, 4, 1, 0, 25, 1, -13, 0, -20, -17, -23, 18, -1, -22, -10, 13, -4, 22, 50, 18, 34, 20, -57, -5, 23, -17, -3, -3, -11, 14, 10, -1, 12, -5, 9, 3, 25, 4, 3, 21, -14, -9, -16, -5, 27, -6, 14, 1, -36, 15, -10, -7, 19, -3, -13, -10, -1, 9, -7, 7, -4, 5, 4, 14, 4, 6, 21, 26, 11, 13, 2, -37, 17, 3, 2, -25, 5, -15, 11, -64, -20, -6, 12, 10, -34, -4, -8, -11, -38, -5, -22, -8, 1, -22, 11, 13, -17, 17, -8, -7, 5, 4, -2, 14, 11, 9, 29, -15, -1, -6, -18, -1, 4, 13, 30, -5, 6, 24, -13, 16, 2, 8, -6, -27, 21, -12, 12, -44, -12, 0, -5, 24, -19, 6, -22, -24, -35, -46, -32, -10, 9, -27, 16, -12, -24, 29, -14, -22, 1, 7, -13, 16, 19, -10, -2, -22, -28, -14, -5, -27, -14, 34, 52, 1, 27, 55, -53, 23, 17, -2, -31, -29, 18, -10, -6, -14, -31, -10, -6, 31, 11, 11, -11, -24, -20, -47, -47, -5, 17, -24, 28, -29, -27, -32, -3, 22, 11, -6, -4, -3, 0, -1, 2, 39, 8, -15, -11, -6, -16, 29, 49, 11, 31, 23, -37, -1, 10, -7, 6, -7, -2, 10, 0, 10, -14, -11, -3, -1, 22, 2, -23, 12, -8, -12, -23, -10, 25, 5, 7, 0, -11, 5, 8, 11, 3, -21, -19, 0, 3, 11, -11, 19, 7, -6, -6, 8, 15, 2, 7, 20, 24, 2, -21, -60, 13, -5, 1, 5, -1, 0, -11, -4, -8, 8, -2, 15, -31, -12, -3, -9, -7, 7, -14, 5, 1, -6, 14, 6, -5, 0, 3, -18, 2, -7, -11, 10, 4, 3, 9, -2, 1, -6, -5, 4, -3, -5, 18, 0, 2, 12, -5, 6, 12, 0, -12, -10, 17, 2, -6, -22, 10, -1, 14, 13, -27, -4, -7, -8, -13, -28, -32, 2, -4, -17, -3, -14, -26, -4, -10, -12, 5, 16, 9, 1, 4, 3, 0, -28, -24, 1, -12, -17, -17, 10, 8, -27, -11, 4, -19, 12, -37, 10, -46, -17, 12, 1, -19, 2, -9, -22, -12, 33, -15, 14, 5, 9, 8, -18, -31, 8, 9, -27, -7, -9, -13, -13, -6, 14, 10, 32, 10, 6, -4, 12, 6, -11, 8, -4, 0, 0, -24, 20, 13, -12, -10, 3, -5, 10, -14, -6, -2, -5, -18, 8, 10, -1, -4, 8, -13, 10, -5, 2, -3, 5, -10, -4, -12, -16, -2, -2, -19, 8, -6, 10, 0, -6, 5, 0, 5, 6, -3, 11, 1, -3, 5, -9, -5, 3, 1, -5, -2, -17, 2, -1, -5, -10, 20, 4),
    (-29, 6, 11, -11, -15, 11, 6, -11, -35, 20, -10, 8, -23, -26, 17, 5, -26, -12, -16, -6, 18, -1, 5, -15, -19, -20, -28, 8, -27, -1, -19, -3, 8, 34, 28, 24, -18, -11, 28, -5, -2, 16, -17, 14, 19, -12, -14, -4, -71, -13, 5, 4, -28, 6, 9, 3, -33, 14, -3, 17, -33, -31, 10, 21, -14, -3, -37, -7, 4, -28, -14, -20, -20, -24, -16, 6, -31, 8, -42, 22, 1, 28, -2, 49, -19, -24, 23, 1, -10, 27, -54, 24, 21, 4, -20, -11, -33, 21, 5, -3, -35, 8, 14, -2, -6, 2, -8, -28, -3, -16, -7, 22, -5, 3, -1, 3, 6, -11, -15, -17, 20, -14, -6, 5, -19, -5, -22, 7, -5, 22, -4, 30, -21, -15, 39, -18, 4, 7, -20, -2, 11, -5, -20, -23, 7, -2, -18, 11, -27, -20, 2, -6, -15, 2, -14, 9, -6, -10, -3, 22, 8, -24, -5, -8, -9, -32, 7, -11, -6, -18, 18, 13, -7, -25, -16, 8, -10, -2, 3, 8, -43, -2, 8, -8, -7, -8, -30, -3, -6, -3, 9, -22, -29, 1, 1, 1, -16, -12, -3, -5, -24, 23, 4, 35, -36, -51, 8, 10, 23, -14, -51, -16, 5, -35, 6, -9, 7, -47, -17, 11, -16, -1, -18, 22, 12, 32, 22, 36, -4, -20, 35, -6, 16, 11, -36, 22, 11, 1, -32, -9, -47, -33, -20, 13, -18, 8, 16, -4, -22, 1, 11, 19, -36, -57, 14, 28, 16, -4, -61, 6, -20, -30, -18, -17, -34, -13, -23, 8, -6, 2, -44, 33, -2, 53, 6, 31, -18, -32, 41, -5, 3, 21, -67, 20, 23, 13, -31, 9, -32, -11, -20, 6, -26, 14, 25, -8, 3, -3, 14, 3, -18, -10, -5, 27, 10, 30, -43, 7, 2, -24, -19, 28, 5, -26, 0, 22, -6, -8, -31, 9, -4, 36, -1, 27, 6, -10, 46, -25, 16, 2, -28, -12, 24, 15, -9, -1, 13, -12, -7, 6, -11, 1, -7, -9, 5, 0, 0, 2, 5, -6, 3, 17, 4, -29, -12, -10, 4, -15, 1, 4, 3, -5, -16, 20, 3, 2, -10, -9, 8, -7, 17, -3, -30, -15, -8, -1, -12, -6, -30, -1, 1, 6, -19, -7, -16, 2, -12, -4, -12, -8, -13, -1, -11, 13, -10, 24, -16, -43, 13, -2, 8, -3, -45, -14, -3, -44, -2, -12, 11, -26, -14, 8, -7, -12, -4, 19, 15, 25, 17, 21, -20, -5, 15, 0, 3, 0, -19, 8, 8, -2, -22, 18, -36, -21, -9, -1, -6, -1, 14, -14, -10, 5, -6, 10, -41, -41, 5, 1, -1, -7, -63, 2, -25, -53, 3, 6, -6, -4, -15, 12, 7, -1, -28, 18, -3, 40, -5, 17, -21, -33, 31, -9, -3, -10, -16, 15, -7, -1, -24, 9, -14, -7, 2, -8, -18, 8, -7, -2, -20, 9, -2, 2, -31, -18, 31, 6, 8, 14, -23, 1, 34, -39, 16, -12, 12, -16, -5, 23, 24, -7, -29, 16, 14, -8, 13, 19, -18, -11, 23, -17, 4, 15, -10, -13, 2, -2, 3, -10, -1, -5, 11, -5, -12, 4, 25, -9, -17, -5, 14, 16, -13, -5, 28, 10, -7, -4, -16, -5, -33, -25, 7, 1, -12, -33, -15, 4, -17, -22, 10, -2, 12, -18, 24, 18, -21, -8, -8, -24, -11, 3, -24, -3, -11, -4, -2, -4, -2, 10, -13, -18, -16, 6, -4, -3, -2, -6, -14, 0, 1, -15, 11, -4, -2, -8, -9, 6, -20, -22, 7, 1, 17, -4, -12, 7, -5, -20, -2, 12, -2, 0, 0, 2, -22, -4, -14, -8, -10, -10, -20, 0, 9, 5, -20, 13, -14, -2, 2, -12, -27, 9, -5, 6, -3, 9, -22, -1, -14, -11, -2, -18, -7, -7, -31, 2, -12, -27, -9, 5, -1, -2, -2, -4, -9, -17, 6, 14, -24, 6, 2, 7, -20, -24, 5, -13, -15, -5, -28, 4, -1, -7, -24, -12, -7, -6, 11, -22, -29, 12, -11, 10, -5, -1, -15, -10, -13, -10, 14, 25, -11, 5, -19, 6, 2, -23, 12, 3, -8, -15, 8, 3, -4, -18, 5, 11, -21, -5, -6, -16, -24, -12, -13, -24, -8, -2, -8, -5, 12, -11, -18, -8, -2, 10, 8, 4, 12, 7, 1, 14, 8, -10, -2, 8, -4, -9, 10, 15, 16, -13, -25, 12, 7, 5, 13, -17, -4, 16, -15, 9, 19, 0, 5, 6, -2, 16, -2, -8, -22, -13, -5, 4, 9, 15, 3, 9, 8, 7, -8, 2, 9),
    (9, -12, -22, 12, -2, -2, 3, -5, 10, 15, 13, -1, 18, -21, 1, -5, -5, -29, -10, 4, 7, -3, 10, 41, -16, -16, -19, -37, -3, -15, 16, -21, -5, -11, 22, -14, 11, 3, 12, 24, 12, 5, -8, -1, -25, 29, 0, -8, -25, -16, -4, 2, -14, 0, 5, -7, -11, 12, -5, 4, 19, -13, -4, 9, -11, -48, 2, -3, 2, 14, -5, 25, -19, -13, -16, -48, 7, -32, 25, 22, -12, -17, 13, -10, 1, 3, 11, 22, -9, 7, 19, 32, -34, 18, -11, -12, -26, -12, -1, -10, -11, 1, -8, -7, -9, 8, -6, -7, 3, -2, 3, 0, -5, -12, -4, 15, -12, 14, -3, 14, -25, -13, -1, -16, -3, -32, 6, 11, -10, -15, 5, -2, 2, 3, 5, 26, -7, 18, 18, 22, -8, 22, -20, -6, 0, -8, 1, -12, -1, 0, 1, -11, 7, -6, -13, -8, 5, -2, 6, 7, -2, 13, -15, 2, -11, 11, -3, -9, -8, -13, -4, -3, -12, -24, -2, 7, -9, -2, 8, -5, -3, -13, 9, 10, 4, 2, 5, 11, 6, 8, 6, 2, -3, -22, -19, 14, 11, -10, 15, 11, 24, -39, -7, -8, 12, -26, 18, -5, 25, -17, 6, -4, -13, -15, 8, 45, 2, -32, -23, -32, 4, 13, 14, 12, -35, 5, 31, -27, 7, 18, -5, 14, 15, -17, -14, -15, -38, 31, 0, 2, 3, -17, -8, 22, -2, 19, 3, 2, 28, -18, -4, -30, 18, -35, -22, 2, 30, -25, 18, -6, -15, 7, 7, 49, 0, -15, -23, -46, 10, 3, 1, 30, -38, -1, 37, -19, 6, 7, 6, 38, 2, -13, 2, 8, -54, 41, -11, -22, -5, -23, 2, 13, -4, 5, -13, 0, 37, -13, 4, -24, 6, -15, -10, -6, 17, -37, 23, -20, -14, 4, 0, 33, -26, -6, 2, -30, -10, -9, -11, 29, -28, -10, 34, -12, -9, -1, 7, 30, 0, 2, 15, 11, -39, 42, -14, -12, -18, -11, -10, 6, 1, -9, 11, -15, 3, -6, 0, -5, 4, -8, -4, 9, -5, -38, 14, 6, -19, 1, -9, 21, 3, -5, 6, -3, -12, 1, -24, 11, -22, -12, 15, -1, -10, -4, 9, 10, 7, 3, 11, 8, -12, 24, -21, 5, 16, -16, -28, -7, 11, 12, 20, 14, 17, -11, -13, -13, 22, 6, 1, 0, 18, -7, 4, -3, 1, -11, -14, 18, -1, -8, 5, -16, 6, 20, -3, 1, -34, -1, 2, -4, 16, 10, 7, 5, 27, -24, -17, -15, -22, 12, -1, -11, 13, -15, -18, 11, -3, 42, 13, 27, 26, -7, -10, -22, 18, -15, -11, 7, 26, -1, 20, 1, -12, -3, 1, 26, 9, 10, -5, -15, -7, 16, 7, 25, -28, 30, 8, -12, 14, 3, 16, 21, 18, -24, -4, -13, -12, 37, -1, -32, 8, -24, -3, 10, -12, 28, 8, 26, 21, -9, -11, -17, 7, 4, -8, 10, 22, -11, 12, -18, -15, -9, 9, 26, 9, 10, 19, -34, 4, 10, -1, 14, -11, 15, -12, -17, 4, -9, -13, 29, 8, -8, 0, -3, 4, 36, 30, -26, 8, -3, 7, 20, -2, 12, -1, 5, 20, -7, 1, -15, 21, 12, 1, 20, -1, -6, -1, -13, 8, -4, -2, 18, 2, -2, 2, -12, 36, 11, 28, 6, -7, -1, 2, -8, -15, 10, -1, 4, 11, -3, -18, -17, -7, 29, 8, -10, 2, 10, -12, 10, 7, 2, -3, -2, 8, -1, -11, 9, 8, 13, 3, 1, 9, -5, -10, 4, 0, -2, 12, 16, -1, -24, 2, -1, 9, 3, 1, 1, -21, -5, 1, -1, 18, 3, 7, 8, 3, -5, -7, -13, -9, -1, 4, 4, 12, 14, -8, 6, 15, 21, 10, 5, 19, -16, 4, -13, -2, 12, 2, 18, 8, 2, -1, -3, -11, 3, 2, 23, -1, 8, -6, 9, -22, 10, -2, 3, -3, 7, 20, -1, 14, -1, 10, 24, -7, -17, -4, -8, -9, 9, 0, -4, -5, -4, 0, 13, -11, 12, 1, 7, 11, -8, -10, -3, -20, 9, 8, -5, 8, -10, 6, -4, 8, -2, 1, 17, -2, -2, -5, -18, -12, 13, 17, -2, -13, 5, 13, -7, 6, 11, 0, 8, -4, -5, -1, -5, -7, -1, 3, -9, 6, -9, -5, 13, -8, 8, 5, 9, 2, -1, 0, 1, 13, -19, -8, 6, 5, -20, 2, 0, -1, 2, 4, 8, -3, 20, 1, -9, 2, 5, 5, 5, -7, 1, 7, 9, -6, 17, 0, 2, 13, 5, 5, -4, -1, 1, -3, -6, -3),
    (-10, -21, 22, 8, -19, -5, 13, 9, -10, -37, 7, 5, 13, -23, -9, 17, -2, 34, 8, -10, 24, 11, 2, 10, -50, 0, -1, -4, 7, -5, 28, -15, 0, -47, 24, -20, -13, 25, -12, 16, 24, -6, 19, -10, -24, 33, -20, -17, -35, -16, 26, -9, -28, -7, 24, 3, -24, -57, -13, 31, 8, -17, -8, 13, 6, 28, 11, -30, 26, 14, -2, 4, -50, -3, -20, -13, -5, -6, 8, 10, 2, -39, 19, -25, -3, 30, 11, 22, 2, -17, 30, 11, -20, 19, -23, -1, -16, -13, 27, -11, -4, -2, 19, 12, 5, -25, -6, 15, 7, -8, -7, -5, -2, 4, 15, -23, 17, 20, -4, -1, -32, 4, -3, -13, -6, -7, 3, 6, 2, -24, 15, -17, 11, 26, 1, 22, -8, -5, 30, 11, -15, 15, -25, -4, -4, 24, 18, -2, 8, -1, 13, 0, -15, -8, -11, -21, 1, 5, -8, -17, -12, 8, 3, -9, 8, 14, -2, -17, 7, 1, -12, -24, -4, 6, -2, -2, 2, -28, -9, -21, 10, 7, -20, 12, -1, -14, 21, 10, -11, 5, -7, -1, -10, -12, 35, 13, -10, -9, 13, -1, -27, -1, 26, 20, 15, -10, -13, 23, -33, 11, 21, -48, 11, 19, -8, 2, -36, -12, -1, 2, -4, -14, 12, -29, -27, -30, 13, 2, -11, 32, -29, 4, 2, 22, 27, 2, -31, -7, -22, -1, -18, 1, 27, -1, -7, -56, 18, -19, -38, -9, 11, 19, 14, -15, -33, 9, -10, 16, 8, -55, 19, 19, -3, 5, -47, 5, -15, -14, -24, -1, 3, -25, -13, -35, 25, -34, -3, 30, -16, -2, -14, 33, 13, 18, -13, 5, -31, 1, -3, -5, 13, -13, 0, -40, 16, -4, -24, 0, 10, 23, 3, -8, -27, -1, -10, 25, 10, -42, 16, 18, -3, -14, -50, 6, -21, 3, -29, -2, -5, -6, -4, -34, 9, -15, -2, 24, 2, 3, -10, 0, 7, 16, -22, 22, -24, -1, -9, 5, 8, -19, 2, -19, 0, -5, -12, -4, 4, -2, 6, 3, -13, -12, -6, -2, 7, -4, 4, 11, -2, -13, -9, -2, -12, -11, -16, -1, -4, -13, 12, -27, -4, -13, 27, 4, -19, 8, -21, -4, 3, -2, -1, -8, -17, 4, -4, -19, 0, 1, -7, -12, 11, 25, -13, 4, 24, 15, 16, 0, -15, 35, -29, 2, 6, -18, 15, 14, -6, 3, -13, -23, 3, -11, 4, 16, 14, -24, -17, -14, 12, -11, -16, 26, -38, -3, 17, 16, 10, -1, -17, -1, -2, -3, 10, -11, 18, 4, -7, -35, 18, -8, -13, 0, 33, 14, 24, 3, -35, 24, -13, 2, 5, -8, 25, 20, -1, 5, -20, -8, 6, -10, 11, 11, 21, -20, -4, -3, 30, -20, -6, 23, -29, -17, 16, 18, 8, -1, 1, -4, 2, 7, -5, -16, 4, -4, 9, -23, 23, 4, -14, -4, 31, 18, 23, 12, -24, 25, -7, 5, 1, -1, 0, 29, 13, 6, -21, 3, 7, -3, 19, 13, 2, -12, -1, -5, -1, -10, 1, 23, -24, -11, 6, -2, -3, 9, -16, 6, -1, 4, -1, -4, -6, -1, 16, -17, 2, 8, -8, -1, 4, -5, 7, -6, -17, 7, -10, 10, 12, 3, 14, 12, -11, 2, 4, 0, 4, -8, -8, 12, 3, -6, 6, -20, -17, -27, 13, 19, -27, 8, 2, -22, 3, -10, 1, 3, -1, 8, 1, 17, -7, 4, -14, -6, 6, 8, 18, -12, 19, 8, 6, 11, -15, 14, -3, 6, 0, -7, 16, 7, 9, -2, -8, -13, 19, -9, 29, 21, 15, -9, 2, 0, 20, -9, 12, 20, 10, 7, 12, 6, 11, -9, 0, 11, 9, -13, 1, -2, -12, 15, -8, -17, -17, 7, 3, -11, 28, 17, 15, 11, -20, 25, -7, 1, 3, -2, 7, 2, 4, -5, -3, 4, -6, 25, 35, 17, 13, -16, 12, 25, 7, 5, 0, 11, 16, -11, 17, 12, 5, 3, 12, 0, 7, 8, 6, -21, -1, -2, 6, -12, -1, -16, -6, -1, 14, 0, 14, 8, -14, 1, 2, 9, 11, -13, -8, 9, -7, 11, -9, 17, 0, -6, 30, 9, -5, -11, 14, 8, -10, -10, -1, -4, -17, -1, 15, -12, -3, 3, -14, -5, 6, 4, -2, -23, 31, 3, -4, -4, 2, -25, -5, -20, -7, -3, 10, -17, 2, 6, -8, -11, 17, -14, 17, 20, -1, 7, -5, 3, -3, -11, 0, -14, 8, -7, 5, 2, 0, -11, -13, 18, -26, -8, 6, -23, 2, -9, 10, -19, -12, 14, -14),
    (11, 3, 14, 7, -24, -14, -5, -4, 17, -14, -50, -12, -10, 11, -21, 34, 11, 28, 34, -12, 8, 21, -11, -23, -23, 11, 38, 22, -6, -20, -37, -20, -5, -12, -1, -16, 19, -8, 3, -23, -20, 7, -3, -3, 14, -25, 3, -15, 30, -15, 30, -17, -24, -25, -17, -23, 25, -19, -50, -23, -13, 24, -34, 36, 2, 28, 33, 8, -3, 5, -39, -17, -14, 18, 40, 34, 16, -21, -63, 10, -14, 1, 9, -47, -5, -4, -15, -3, -9, 0, -55, -7, 19, -14, 4, -32, -7, -2, 15, -22, -8, -27, -24, -23, 3, -12, -54, 13, -14, 2, -32, 29, 22, -11, 25, -4, 5, 10, -28, -13, 3, 7, 31, 24, 2, -17, -63, 14, -4, 23, 5, -23, -12, -11, 3, 23, -6, 6, -52, 1, 12, -9, 12, -40, -7, 8, -9, -13, -4, -23, -7, -9, -3, -3, -23, 10, 2, -7, -9, 21, 10, -21, 5, -8, 17, -12, -13, 11, 5, -13, 25, 6, -19, -7, -18, 12, -4, 20, -1, -8, -26, -3, -2, 19, -12, -2, -27, 1, 15, -14, 6, -15, 21, -15, 12, 7, -1, 4, -11, 1, 10, -24, -14, 27, -9, 30, -1, 40, 32, 22, 51, 39, -18, -1, -23, -4, -31, 24, 62, 19, 6, -2, -15, -24, -17, -42, -10, -11, 5, -4, -9, 3, -3, -7, 11, -8, 18, 1, -17, -39, 28, -13, 15, 5, 3, 11, -1, -13, 13, -8, -37, 0, 2, 36, -56, 35, 15, 39, 39, 29, -13, -5, -22, 14, -41, 19, 57, 21, 36, -4, -45, -18, 1, -13, -6, -34, -4, -1, -27, 12, -4, -15, -3, -33, 37, 13, -17, -43, 17, -27, 17, -2, 5, -13, -13, -17, 14, -5, -28, 8, -5, 5, -42, 31, 14, 47, 27, -1, -6, -3, -33, 14, -28, 4, 30, 6, 16, 4, -51, 6, -2, 15, 9, -16, -6, -12, -5, 22, -1, -10, -21, -24, 33, 16, 10, -29, -10, -1, -8, -6, 5, -4, -12, -12, 14, 9, -8, -4, 0, 6, -27, 5, 18, 18, 5, 1, -6, -6, -10, 0, 1, 3, 24, 15, 4, 5, -9, 18, 5, 12, 8, 1, -18, -16, 23, 7, -8, 6, -35, 3, 3, -1, -4, -17, 1, -18, 22, 5, 4, 4, -6, -17, 1, -17, -37, 28, 0, 31, 11, 15, 24, 4, 33, 18, -12, -22, -16, 4, -49, 20, 17, 17, -20, -19, -2, -14, 1, -43, 9, 10, -4, -11, 2, 22, -32, -24, 11, -7, 3, 8, -18, 5, 6, -10, 23, 0, 15, 20, -2, -15, 13, -14, -44, 14, 4, 47, 28, 23, 21, 14, 30, 11, -8, -12, -6, 0, -43, 27, 17, 16, -31, -19, -8, -14, -1, -43, -17, 6, 5, -26, -7, 28, -23, -39, 15, -41, 6, 27, -17, -21, 10, -3, 7, -9, 6, 4, 0, 9, 10, 10, -20, 4, -14, 8, 11, -2, 24, 19, 14, -1, -14, -17, 12, 2, 1, 16, -12, 0, -1, -1, -4, 0, 2, -14, -4, 9, -1, -22, -12, 31, -7, -31, 3, -22, 3, 18, 1, -12, -4, 0, -9, 1, 3, 9, -4, -5, 8, 3, 5, 1, 0, 18, 5, 0, 10, 16, 5, 3, -13, -15, -6, 5, -8, -1, 10, 6, 10, 7, 6, 8, 7, -14, 1, -10, 5, 1, -6, -1, 11, 5, -24, -11, -14, 3, 10, -6, -6, -21, 12, -19, 13, 8, 8, -7, -4, 8, -12, 20, -7, -13, 10, 5, -10, 10, 10, 0, -32, -19, -7, -3, -39, 13, 18, 8, -44, -25, -4, -7, 12, -10, 0, -4, -20, -30, -17, -4, -19, -14, 1, -18, -12, 1, -25, -9, 0, -29, 10, -20, 5, 17, 36, -8, -11, 4, -31, 9, -14, -2, 9, -6, 14, 3, -4, -3, -32, -16, 8, -11, -28, -17, 21, -1, -21, -30, -5, -11, -8, -25, -2, 6, -6, -20, -8, 18, -27, -28, 16, -1, -17, 14, -28, 9, 6, 11, 11, 2, -10, 5, 11, -5, 1, 4, -19, -10, -5, 10, 3, 1, 11, 3, -6, -5, 9, 5, 2, 7, 8, 5, 8, -8, -36, -10, 8, -1, -6, 2, -10, -5, -8, 11, -18, -2, -16, -8, -1, -3, -12, 2, -9, 2, 9, -7, 3, -6, -8, -7, -10, 10, -6, 7, -8, -3, -11, 16, 0, 9, 3, -22, 11, -11, -5, 3, 7, -2, -4, -17, 10, -2, -11, 0, -9, 8, 4, 0, -7, 4, -3, 1, -10, -8, 10, 13, -12, -8, 0, 7, -1, -7, 2),
    (-4, 18, 4, -17, 4, -24, 1, -8, -5, -11, 29, 3, -7, 5, -31, -1, -8, 9, 6, 16, 13, 10, 6, -15, 19, 5, 1, -5, 7, 11, -5, -15, -16, 29, -1, 5, -4, 17, 1, 15, -6, -5, -6, -11, 13, -19, 1, -11, -7, 39, -3, -16, 13, -47, -1, -11, 5, 2, 30, 19, -9, 13, -37, 0, -2, 12, 13, 15, 28, 4, 6, -21, 35, -8, 10, 10, 8, 46, 1, -35, -3, 38, -14, 0, -18, 20, -12, 10, -1, -32, -31, -48, 8, -20, 16, -28, 9, 13, -16, 0, 29, -43, -7, -4, 10, 3, 30, 41, -3, 9, -31, 34, 16, -28, 23, -15, 24, -7, 8, -13, 34, 3, 11, -18, 17, 55, 7, -20, 8, 39, -15, -23, -11, 9, -21, -28, -3, -39, -52, -41, -1, -39, 24, -19, 3, -3, -15, 9, 7, -22, 2, 9, 16, -4, 25, 16, 2, 6, -33, 21, 11, -9, 4, -18, 22, -7, -4, 13, 16, 1, 13, -3, 5, 24, -13, -4, 16, 15, -22, -26, -26, 18, -19, -17, 7, -23, -22, -35, -12, -21, 3, 10, -17, 18, 23, -6, 8, -24, 8, -16, -12, -10, 25, -3, 8, 0, -12, 4, -10, 9, 8, -14, 14, 10, 12, -20, 2, -1, -10, 6, 22, -1, 1, -60, 9, 3, -9, 2, 6, 20, -22, -4, -12, -3, -6, 0, 6, 2, 0, -15, -28, 26, 12, -20, 11, -54, -6, -22, -15, 5, 22, 12, 5, 9, -34, -1, -13, 26, -6, -15, 15, 7, 20, -40, 22, 3, 8, -7, 34, 16, 16, -61, 13, 34, -19, 12, -1, 32, -33, -16, -18, -7, -12, -42, 15, -14, -4, -8, -17, 23, 9, -8, 0, -41, -11, 0, -24, 22, 28, 27, -3, 16, -19, 6, -5, 9, 6, 20, 21, 1, 18, -6, 39, -2, 6, -20, 38, 5, 18, -40, 17, 20, -55, -2, -12, 32, -48, -22, -4, -26, -28, -29, -2, -28, 23, 5, -9, 32, -23, 24, -5, 4, -19, 0, -9, 19, 28, -7, 1, 14, -9, 11, -5, 3, -4, 1, 4, 6, 2, 8, 10, 1, -1, -20, 47, -1, 13, -14, -6, 10, -12, -7, -4, 8, -31, -35, 10, 1, -20, -12, -14, -12, 35, -3, -9, 12, 7, -10, -13, -24, 13, 6, -1, -3, 17, 3, 10, -6, -8, 8, -11, 19, 12, -1, 15, 25, 4, -7, -1, 15, 3, -20, 2, 7, 19, -22, 1, -16, 1, -14, -4, 25, -18, 3, 0, 3, -10, -11, -21, 13, 0, 10, 1, 22, 2, -11, -8, -33, -11, -10, 0, 9, 19, 11, 9, -2, 11, 11, -17, 31, -6, -16, 16, 23, 2, -8, 13, 0, -4, -13, 21, -3, 18, -25, 2, -4, 13, -17, -11, 14, -21, -14, 0, 3, -10, -11, -15, 0, -6, 1, -23, 2, -7, -5, -13, -23, -10, -3, -15, 3, 15, 25, 15, 4, 14, 12, -21, 13, -10, 9, -11, 10, 2, 0, -15, -12, -8, -15, 17, 1, 16, -22, -2, 12, 9, 4, 3, 13, -10, -32, 1, 10, -23, 4, -15, -18, -14, 1, -14, 4, -4, 7, -16, 4, -9, -2, -5, 2, -6, -17, -1, 4, 11, -21, -3, 5, -17, -5, -10, 10, 3, -2, -13, 6, 4, -9, 8, -7, 1, -11, -4, -4, 6, -1, 5, 3, -1, -9, 2, 0, 7, 2, 3, -5, 19, 10, 2, -1, -8, -10, 1, -11, 11, 0, 2, 8, 22, -3, 8, -5, -12, 10, -10, 2, -4, -8, 19, 7, 7, -6, 2, -5, 2, -5, -10, 12, 5, -12, -1, -9, 3, -6, 8, 26, -7, 4, 5, 3, 3, -12, -14, 15, -1, -7, -1, 7, 12, 5, 3, -15, -3, -18, -6, 14, 12, -2, 16, -2, -19, 12, -16, 15, 12, 0, 14, 4, 13, -5, 7, 24, -1, -9, -17, 18, 8, -9, 11, -7, 6, -9, 8, 21, -17, -14, 11, 5, 11, -17, -2, 3, 8, 3, -8, -16, -1, 12, 16, -21, -3, -12, -2, -4, 8, -1, 15, 13, 0, -12, -26, -10, 12, 2, -11, -6, -7, -5, -7, 4, 15, -7, -1, 2, -2, -2, -1, -12, 11, -18, 0, 9, -16, 2, -3, -9, 3, -3, -14, -1, 2, 12, -10, -3, -8, 1, -5, -14, -3, -9, -9, 6, -8, -3, -8, -7, -4, -17, -5, -15, 11, 6, -23, -16, 6, -16, -7, -13, 0, -7, -4, 14, -7, -11, 6, -19, 3, -20, -3, 0, 1, 6, -14, -10, -3, -1, -17, -8, -11, 10, -3),
    (-15, 7, -2, -41, 11, -6, -28, -21, -13, 20, 4, -12, -14, 19, -13, 5, -25, -18, 22, -11, 9, -12, -3, -7, 22, 12, 7, -24, -8, -7, -39, 29, -17, 30, -6, 10, -16, -14, 28, -13, -9, 5, -22, 2, 15, -63, 4, -16, -44, 24, 4, -35, 9, -13, -50, -44, 25, 20, 8, 6, -21, 26, -31, -5, -9, -2, 27, -16, 8, -19, 14, -22, 23, 2, 10, -40, 2, -12, -46, 17, -42, 25, -29, 18, -16, -10, 35, -30, -28, 1, -49, -3, 4, -69, 8, -40, -24, 23, 1, -5, -47, -1, -24, -23, 9, 5, -11, 6, -20, 21, -14, -22, -12, 32, 12, -18, -8, -7, -3, -16, 25, -9, 4, -42, 8, -10, -18, -7, -23, 16, -6, 19, -30, -7, 10, -7, -17, 2, -32, -10, -4, -29, 16, -50, -4, 0, -7, -7, -22, -15, -2, -8, 6, 3, -4, -5, -18, -3, -1, 22, -19, -3, -4, -7, -11, -18, 3, 8, 11, -18, -8, 1, -4, -6, -20, -11, 3, -2, 1, -2, -48, 7, 1, -10, -11, -13, -8, -25, -9, -26, 3, -36, 10, 4, -20, 7, -1, 14, -45, -39, 29, 19, 8, -28, -6, 15, -9, -21, -10, -9, 23, 14, -18, -15, 17, 12, 13, 7, 18, -14, -1, -1, -33, 14, -5, 17, -16, 11, 13, -25, 22, -20, -19, 9, -2, 6, 14, -35, 2, 7, 32, 10, -5, -9, 17, 19, -69, -39, 32, 15, 9, -18, 2, 19, -10, -14, -9, 15, 25, -2, -9, -10, 22, 3, 17, 9, 26, -35, 9, 1, -23, 18, -28, 23, -30, 27, 18, 7, 31, -28, -38, 12, -3, 4, 7, -51, 12, -25, 24, 10, 7, 17, 3, -1, -41, -10, 22, 5, 1, -32, -13, 25, -6, -34, -12, -15, 11, -4, -10, -7, 24, -2, 20, -2, 13, -42, 7, -10, -4, 0, -26, 20, 0, 14, 7, 7, 13, -11, -26, 2, -16, -5, -5, -46, 19, -16, 4, 17, 2, 10, 3, 9, -2, -1, 12, -11, 4, -22, -6, 6, 6, -10, -7, -14, 6, -3, -8, -10, 3, 0, -16, -3, -1, -2, -4, -8, 5, -14, -8, 10, -2, 16, -23, 7, -5, -3, -9, -10, 1, -9, -12, -4, 4, 1, 7, 2, -15, 24, 8, 7, -39, 4, 10, 11, 5, -38, -18, 26, -7, -42, -33, -2, 34, 1, -16, -15, 12, 5, 10, 16, -6, -35, 0, 7, 3, 23, -2, -1, -17, 1, 14, -22, -6, -17, 0, 7, -6, 17, 23, -11, 19, -6, 25, 16, -16, 18, 9, 21, -33, 3, 14, -2, 7, -17, -16, 25, 16, -30, -15, 15, 13, 4, 8, -8, 4, 11, 5, 16, -11, -34, 4, 2, 2, 15, -33, -2, -6, 27, 21, -3, 12, -26, 4, 1, -15, 6, 30, -25, 23, -22, 22, 1, -19, 14, 8, 5, -1, 10, 3, 9, 15, -15, -13, 25, 12, -18, -18, -14, 4, -2, -20, -4, 5, 24, 4, 11, -6, -31, -4, 4, -13, 1, -22, -8, 7, -13, 19, -11, -5, -12, 7, -1, -21, 7, 3, -21, 18, -4, -7, 0, -14, -9, 5, 5, -5, 11, 0, 2, 2, -7, -21, 17, 1, -13, 0, -19, -6, 0, -16, -5, -12, 7, -9, 11, 4, -5, 0, 12, -1, -10, -4, -4, 6, -4, 6, -5, -9, -12, -1, -5, 0, -6, 0, -5, -27, 0, -1, 0, -16, 9, 17, 3, -17, -3, -6, -6, 16, -39, -23, 3, -21, -15, -18, -17, 14, -3, -13, 5, 8, 4, 3, 10, 0, -11, 4, 2, -6, 16, -25, -23, -2, -21, 1, -13, -29, -23, 10, -7, -28, 7, 5, 0, 14, 7, 5, 1, -1, 17, 13, 7, -9, -5, 3, -10, -1, -40, -5, 9, -7, -13, -25, -10, -3, -6, -5, -17, 4, -3, -5, 8, -10, -22, -4, 2, -9, 8, -7, -18, -11, 3, 13, -3, -24, -16, -5, 0, -22, -13, 13, -7, 14, -17, 2, -18, 5, 4, 4, -2, 5, 4, 21, 2, -12, -10, -16, 3, -8, 7, -7, -14, 14, 1, -19, -4, -1, 4, -8, -9, 3, -6, -18, 3, 2, 5, -11, 2, 3, 4, 30, 4, -5, -5, 4, -5, 0, 0, -11, 7, 3, 15, 6, -18, -1, -7, 0, -10, 7, -3, -2, -9, -1, -7, 3, 24, 6, -11, -8, 3, 23, 4, -10, -9, 2, 8, -3, 4, 6, -6, 22, 14, 4, 0, 14, -2, 14, 0, -4, -9, -7, -7, 5, 4, 11, 9, -8, 12, 23, 12, -6),
    (30, -4, -15, 16, -26, 23, -19, 29, 7, -15, 20, 18, 7, 10, 10, 40, 23, 11, -20, 0, -3, -52, 16, 21, -4, 4, 20, 9, -10, 27, 18, 1, 11, -9, 11, -15, -12, 1, 8, -2, 26, -9, -4, -7, -12, 12, -19, 23, 30, -42, -16, 25, -25, 34, -10, 33, -15, -1, -6, 33, -13, 3, 23, 32, 17, -19, -31, 29, -21, -41, 3, 14, -23, -13, 20, 33, 5, 11, 8, -12, 28, -17, -7, -4, -19, 6, -9, -11, 40, -9, 32, -7, -11, -4, -14, 28, 27, -43, -17, 20, -14, 16, 2, 30, -25, -4, -18, 22, -19, -1, 18, 19, -3, 7, -24, 28, 4, -25, 5, 1, -30, -3, 12, 23, 14, 2, 8, 1, 5, -23, -10, 9, 0, 7, 4, -14, 15, -5, 26, 10, 4, -2, 2, 26, 13, -14, -1, -9, 5, -2, 7, 8, -3, 3, -12, 1, -8, 0, -2, -1, 7, -13, -13, 6, -8, -6, 6, 4, -13, 15, 1, 4, -15, -7, 10, -11, 2, 0, 0, -1, 5, -9, -8, -4, 8, 6, 17, 13, 9, 4, 12, 8, -4, -11, -32, 11, -20, 9, -5, 31, -18, -14, -24, 7, -17, -5, 19, 36, 26, -8, -39, 7, -20, -27, -52, 10, -9, -5, -12, 21, -26, -9, 17, 6, 20, -13, 13, -4, -17, 3, 10, -10, 23, -30, 13, 16, -34, -4, -25, -1, -5, -36, -34, 6, -32, 34, -8, 43, -29, -28, -21, 1, -11, 15, 54, 26, -3, -31, -45, 22, -9, -33, -46, -6, -26, -16, -13, 34, 10, -19, 16, 9, 20, -38, 9, -5, -15, -6, 3, -2, 30, -21, 28, 13, -30, 4, -30, 14, -1, -42, -31, -3, -19, 23, 7, 27, -13, -3, -14, 2, -11, -2, 32, 14, 7, -6, -42, 26, 7, -33, -20, -9, -14, -4, -13, 41, 4, -20, 5, 13, 2, -26, 5, 8, -16, -7, 12, -18, 29, -8, 31, 5, -10, -2, -8, 20, 11, -8, -3, -5, -5, 0, 21, 9, 2, -6, -10, 16, 10, 0, 12, 18, 5, 17, -14, 12, -1, -8, 5, 3, 21, 2, -10, 20, -13, -8, 1, 4, 11, 0, 11, -3, 3, -14, 8, -3, 5, 6, 20, 12, 9, 2, -29, 18, -12, -2, -17, -41, -8, -2, 18, -1, -23, -3, -33, 18, -14, -48, 2, 18, 16, 1, -46, 7, -1, -32, -22, -2, 4, -29, -10, 7, 15, -17, -23, -11, 7, 8, 13, 14, -25, -18, 18, -6, -16, -9, 5, 9, -21, 2, -18, -14, -11, -18, -4, -38, -1, -17, 19, 10, -7, -2, -29, 11, -29, -3, 6, 11, 14, -18, -36, 19, -14, -44, -15, -21, -5, -31, 11, 21, 8, -17, -17, -11, 23, -20, 15, 15, -5, -37, 12, 14, -23, -10, 31, 17, -45, -2, -11, -2, -1, -2, 3, -24, 4, -3, -3, 20, -9, 16, -14, 18, -30, -11, -9, -5, 26, 5, -29, 12, 15, -25, 0, -21, 37, -20, -2, 28, -5, 1, 2, 6, 16, -21, -5, 11, -7, -14, -3, 4, -12, 12, 23, 1, -20, 5, 5, 6, 3, -13, -1, 9, -1, -4, 21, -8, -25, -1, 20, 19, -9, -2, 15, -1, 16, 7, -2, 7, 6, -8, -7, 11, 16, -6, -17, 10, -13, 8, -13, 9, -1, -2, 1, 1, 10, 0, 9, 10, -2, -10, 5, 7, -2, 5, -5, 3, -14, -5, 3, -25, -16, -17, -15, 10, -13, 6, -18, 25, -19, -23, 3, -4, -5, -9, -20, 4, -4, -21, -9, -8, -13, -24, -6, 13, 6, -31, -2, -5, 23, 26, -3, 16, -37, -13, 14, -14, -17, -10, 8, 10, -8, 8, -27, -5, -12, 8, 12, -22, -18, 4, 6, 5, -18, -2, -23, 25, -24, -1, 14, -7, 13, 4, -25, 0, 29, -24, -5, -11, 3, -9, 1, 24, 6, -23, -4, -1, 24, -14, 19, 15, -33, -33, 19, 0, -1, -13, -11, 25, 9, -2, -22, -7, -3, 34, 2, -29, -11, 7, 3, 18, 0, -8, -12, 8, -18, -15, 21, 1, 25, 14, -36, -4, 21, -8, 5, -5, 22, -19, 0, 7, -2, -13, 0, -1, 10, -11, 2, 2, -34, -5, -13, 2, -20, 11, -3, -2, 9, 24, -11, -21, 3, -4, -3, 0, -6, 8, 7, 9, -14, -8, -4, -7, -12, 0, -9, 31, -5, -7, -22, 16, 9, -10, 8, 5, -6, -7, 8, -14, 1, -4, 10, 1, -2, 11, -3, 3, -19, 10, -4, -7, 2, 6, 13, -13, 10, -3, -5, 1, 2),
    (-27, 25, 10, 2, 8, -1, 12, -3, -22, -5, -23, -2, 3, -5, 0, -22, 12, -17, -8, -1, 5, 18, 3, -24, 8, 19, -27, 2, 12, -10, 2, -2, 11, -5, -2, -7, 16, 4, -12, 3, -14, 5, -4, 6, 10, -2, 17, 15, -22, 29, 8, 9, 1, 15, 13, 11, -20, 4, -11, -15, -14, 2, 9, -24, 16, -6, -5, -4, 24, 13, -5, -4, 16, 22, -18, -9, -6, 6, 9, 19, 20, -14, 4, -9, 29, -6, -22, -10, -8, 7, 6, -16, 2, 6, 12, 17, 2, 23, 9, 14, 6, 10, 4, 8, 10, 7, -2, -18, -14, -2, 7, -21, 12, 15, -1, -3, 10, 11, 4, 1, 19, 13, -5, -2, -5, 18, 13, 1, 20, -12, 5, 2, 19, -11, -21, 2, 3, 3, 13, -7, 3, -3, 12, 11, -4, 16, 1, 11, 11, 17, 0, 6, -1, 0, 4, -14, -5, 0, -2, -13, 6, 13, 4, -10, -2, 15, 0, 1, -5, 20, -3, 16, 3, 5, 8, -7, -7, -12, -5, 13, 1, -5, 1, 10, 8, 6, 9, 7, 2, -2, -3, 12, -16, 37, 23, -3, 3, -14, 17, 7, -24, 22, -17, -24, -2, -12, -3, -12, 11, -2, -8, -6, 23, 8, 13, -24, -1, 17, -36, -12, -4, 9, -16, 9, 34, 1, 7, -16, 18, -2, -16, -4, -4, -16, -20, -9, -7, 1, 2, -8, -26, 35, 13, -12, -12, -16, 19, 9, -16, 8, -19, -22, -10, -13, -1, -10, 5, -1, 2, -54, 27, 1, -6, -23, 2, 20, -50, -6, -26, 9, -6, 17, 37, -1, 1, -18, 21, -3, -6, -7, -9, -33, -28, -14, 4, -1, -2, 5, -7, 33, 4, -11, 2, -13, 23, 10, 3, 1, -7, -20, -16, 3, 4, -18, -1, -6, 15, -34, 27, -1, -10, 1, 12, 3, -25, 10, -16, 6, 5, -3, 25, 3, 15, -8, 9, 4, -19, -4, -7, -22, -13, -8, 1, -8, -11, 5, 17, 7, -3, -5, 10, -4, -7, 2, 3, -4, 13, -13, -4, 9, -9, 0, 4, 2, 16, -9, 4, 7, 1, 2, -13, 6, -9, -3, -7, 6, -10, 0, -3, 3, 9, 3, -3, -3, -4, -12, 5, 0, -8, -2, -3, -9, -1, 6, -14, 23, 26, 3, 11, 2, 21, 1, 5, 7, 2, -23, 8, -22, 12, -28, 8, 8, -21, 0, 14, -2, 9, -13, 14, 11, -18, 0, 0, 2, 3, 12, 29, 10, -19, -26, 6, 3, -13, 6, -4, 6, -17, -10, 5, 9, 9, 29, -17, 34, 23, 2, 0, 8, 10, -8, 0, -5, -9, -25, -6, -35, 5, -24, 1, 13, -9, -31, 8, -5, 4, 0, 15, 24, -42, -8, -14, 6, -5, 23, 35, 11, -26, -25, 8, 0, -10, -1, -4, 1, -28, -1, 3, 9, -1, 18, -5, 38, 11, -3, 4, 12, 11, -29, 6, -18, -12, -21, -8, -18, 1, -25, -6, -9, 2, -4, 13, 2, -5, 7, -15, 3, -21, -3, -14, 14, -1, 8, 22, -11, -17, -1, 8, -4, 12, 3, -13, 4, -19, 6, 15, -30, -2, 11, 0, 18, -7, -8, 5, 22, 4, -9, -2, 0, 5, -15, -16, 4, -8, -14, 5, -8, 12, 1, -11, -2, 2, 6, 13, 6, -10, -4, -42, 3, -3, -5, -11, 15, -8, -2, 9, 2, 28, -13, -15, 12, -1, 9, 19, -2, -13, 5, 0, 4, 10, 3, 4, 9, -2, -2, 0, 14, 2, -16, 14, -11, -8, -15, 0, 4, -9, 9, 12, 2, -7, -11, 22, 6, -13, 2, 14, 4, 10, 1, 12, 17, -1, -14, 6, -5, -2, 7, 12, 21, -2, 3, -5, 3, 20, -3, 7, 29, 10, -4, 0, 8, 8, 10, -1, 13, 8, -21, 12, 1, 3, -34, -7, -2, 17, -14, -5, 15, -4, -8, 9, -20, -16, 9, -4, -2, 10, 13, 4, 12, 1, -10, 10, 1, -15, 3, 15, 21, -1, -7, 7, -1, 6, 19, 0, 18, 5, -2, 22, 6, -6, 14, -4, 11, 4, 1, -5, 2, 2, -4, -7, -15, 6, 16, -12, 2, -8, 11, -26, -4, -2, -9, -5, 5, 2, 1, 2, -9, 13, 18, 9, 3, 12, -4, -8, 17, -1, 16, 10, -17, 2, 16, -13, 8, 5, -10, 1, 6, 16, -11, -5, 17, -8, 16, -17, 3, -9, 2, 1, 18, -15, 3, -1, -16, -7, -7, -4, -4, -17, 5, -5, 14, -12, -3, -11, 16, -15, 1, 18, -7, 10, -11, 2, 14, -15, 8, -17, -2, 5, -11, 6),
    (20, 3, -11, -8, 21, 17, 8, 14, 22, -12, -8, -8, 0, 16, 10, -40, 5, 20, -17, 21, -26, 19, -6, -18, 25, 8, 7, 17, 4, -10, -4, -9, 4, 4, -25, 2, 13, -25, -20, -26, -15, 7, 9, -4, 5, 3, 9, 27, 26, 7, 3, 9, 35, 18, 22, 17, 10, 12, 8, -20, 3, 0, 21, -49, 13, 36, -27, 26, -12, 4, 1, -17, 25, -4, -1, 20, 4, -6, 12, -30, 10, -17, -26, 15, 21, -23, -37, -31, 1, 6, 14, -14, -7, 4, 35, 32, 25, -2, 2, 16, 25, 12, 16, 20, -4, 6, 1, -8, -5, -8, 16, -52, -5, 22, -33, 16, -13, 0, 6, -17, 15, 12, -15, 6, 14, 10, 23, -20, 13, -18, -9, 8, 24, -7, -10, -16, 9, 1, 18, -4, -2, -2, 17, 21, -3, 8, 2, 8, 6, 18, 0, 12, 11, -5, 4, 1, -4, 7, 11, -21, -8, 16, -4, 5, -9, 23, -5, 2, 7, 6, -5, 1, 13, 8, 16, 2, 10, -12, -8, 2, 22, 6, -18, -3, 4, 2, 18, 11, -7, 20, 7, 20, 13, -16, 9, -14, 14, 3, 7, 11, 16, -9, -38, 21, -4, 35, -11, -1, -20, 9, -18, 32, -11, 21, -23, -18, 2, 24, 30, 21, 13, -15, 0, -31, -7, -7, -35, 16, 17, -20, -18, -24, -8, -1, 17, 0, 9, 14, 7, -6, 6, -6, 6, -33, 17, -11, 20, 26, -2, -6, -35, 12, -2, 31, 16, -13, 7, 19, -28, 53, -1, 5, -12, -30, 6, 1, 23, 17, 27, -13, 21, -51, 9, -40, -51, 21, 11, -34, -36, -22, -5, -48, 10, 4, 11, 7, 28, 0, 11, -12, -4, -42, 1, -7, 29, 29, -10, -1, -23, 15, -5, 3, 14, -21, -4, 21, -16, 34, 2, -12, -6, 3, 7, -8, -23, 18, 4, 6, 10, -34, 11, -21, -19, 8, 12, -30, -16, -19, 10, -24, 9, 1, 11, 1, 19, 12, 2, -15, 0, -18, 14, 5, 8, 22, 3, -11, 2, 3, 8, -5, 4, -6, 3, 18, -6, 8, -14, -10, 2, -5, -7, 4, -29, 8, -1, 3, 8, -11, 1, -1, -19, -4, 7, -3, 5, -7, 13, -7, 11, 4, -10, 5, 4, 8, 1, -26, 24, -18, 3, -7, 15, 13, 2, -18, -31, 24, -21, 9, 11, 2, -17, -10, -34, 15, -13, 14, 1, -17, -14, -13, 13, 17, -2, -43, -6, -26, 6, -23, -5, 22, 11, -22, 13, 2, -33, -18, 13, -4, -9, 16, -6, -6, 3, -20, 27, -19, 13, -16, 11, -9, -14, -8, -47, 16, -15, 31, 27, 5, 12, 10, -10, 21, 12, -1, 1, -18, -27, -18, 34, 11, 4, -26, -5, -45, 15, -46, -36, 37, 8, -39, 5, 10, -35, -34, 21, -18, -53, 17, -14, 14, 4, -11, 19, -16, 14, -1, 14, 5, -22, 4, -27, 18, -31, 3, 24, 10, 9, 2, -25, 14, -1, -25, -1, -16, -3, -11, 9, 20, -21, -4, -8, -25, 12, -22, -25, 7, 1, -26, 0, 18, -28, -23, 16, -14, 5, 8, -9, -2, 5, -7, 8, -6, -8, -13, 9, -22, -3, -5, -20, -13, -22, 8, -8, 1, 14, 11, 0, -8, -13, -11, -3, 5, -7, 3, 15, 6, -6, -18, 5, 8, -3, 1, -13, -5, 11, -14, -2, 7, 2, -18, 1, 6, 5, -11, -4, -5, -12, -22, 0, -28, -10, -9, 8, 21, -17, 1, -9, 27, 7, -9, 18, 2, -8, 9, -15, 7, -12, -28, -11, -21, -28, -6, 8, -6, -38, -25, -7, -17, 14, -11, -5, 17, -25, -28, 14, -10, -25, -5, 17, -8, -17, 10, -23, 6, -25, -38, 19, -18, -14, -13, 13, 5, -20, 3, -29, 29, -8, 4, 6, 1, 18, 21, -10, 4, 7, -24, -1, -15, -15, -16, 15, 5, -4, -29, -14, -15, 10, -14, -12, 7, -22, -22, 16, 22, -13, -6, 29, 8, -7, 13, -31, 14, -2, 5, 18, -19, -19, -2, 6, 1, -7, 6, -12, 9, -14, -4, -5, -3, 15, 8, -15, -1, 5, 0, -3, -12, 2, 7, -3, 2, -5, -17, -15, -9, 1, -15, -4, -2, -34, -7, 21, 7, -21, 2, -4, -2, -19, 9, -9, -1, 14, -11, 19, -8, -10, -8, 9, -4, -7, -12, 8, -11, -12, 3, -8, -11, -11, 1, -10, 2, -7, -4, -10, -6, -17, -15, -6, -7, -23, -10, 1, -4, -19, 8, -13, -1, 14, -15, 3, -1, -8, -4, 8, 4, -18, 0, -6, -2, -2)
  );
  ----------------
END PACKAGE CNN_Data_Package;
